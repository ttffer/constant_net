`timescale 1ns / 1ps
module tb;
parameter DATAWIDTH =64;
reg rst,clk;
reg [7:0]  img0;reg [7:0]  img1;reg [7:0]  img2;reg [7:0]  img3;reg [7:0]  img4;reg [7:0]  img5;reg [7:0]  img6;reg [7:0]  img7;reg [7:0]  img8;reg [7:0]  img9;reg [7:0]  img10;reg [7:0]  img11;reg [7:0]  img12;reg [7:0]  img13;reg [7:0]  img14;reg [7:0]  img15;reg [7:0]  img16;reg [7:0]  img17;reg [7:0]  img18;reg [7:0]  img19;reg [7:0]  img20;reg [7:0]  img21;reg [7:0]  img22;reg [7:0]  img23;reg [7:0]  img24;reg [7:0]  img25;reg [7:0]  img26;reg [7:0]  img27;reg [7:0]  img28;reg [7:0]  img29;reg [7:0]  img30;reg [7:0]  img31;reg [7:0]  img32;reg [7:0]  img33;reg [7:0]  img34;reg [7:0]  img35;reg [7:0]  img36;reg [7:0]  img37;reg [7:0]  img38;reg [7:0]  img39;reg [7:0]  img40;reg [7:0]  img41;reg [7:0]  img42;reg [7:0]  img43;reg [7:0]  img44;reg [7:0]  img45;reg [7:0]  img46;reg [7:0]  img47;reg [7:0]  img48;reg [7:0]  img49;reg [7:0]  img50;reg [7:0]  img51;reg [7:0]  img52;reg [7:0]  img53;reg [7:0]  img54;reg [7:0]  img55;reg [7:0]  img56;reg [7:0]  img57;reg [7:0]  img58;reg [7:0]  img59;reg [7:0]  img60;reg [7:0]  img61;reg [7:0]  img62;reg [7:0]  img63;reg [7:0]  img64;reg [7:0]  img65;reg [7:0]  img66;reg [7:0]  img67;reg [7:0]  img68;reg [7:0]  img69;reg [7:0]  img70;reg [7:0]  img71;reg [7:0]  img72;reg [7:0]  img73;reg [7:0]  img74;reg [7:0]  img75;reg [7:0]  img76;reg [7:0]  img77;reg [7:0]  img78;reg [7:0]  img79;reg [7:0]  img80;reg [7:0]  img81;reg [7:0]  img82;reg [7:0]  img83;reg [7:0]  img84;reg [7:0]  img85;reg [7:0]  img86;reg [7:0]  img87;reg [7:0]  img88;reg [7:0]  img89;reg [7:0]  img90;reg [7:0]  img91;reg [7:0]  img92;reg [7:0]  img93;reg [7:0]  img94;reg [7:0]  img95;reg [7:0]  img96;reg [7:0]  img97;reg [7:0]  img98;reg [7:0]  img99;reg [7:0]  img100;reg [7:0]  img101;reg [7:0]  img102;reg [7:0]  img103;reg [7:0]  img104;reg [7:0]  img105;reg [7:0]  img106;reg [7:0]  img107;reg [7:0]  img108;reg [7:0]  img109;reg [7:0]  img110;reg [7:0]  img111;reg [7:0]  img112;reg [7:0]  img113;reg [7:0]  img114;reg [7:0]  img115;reg [7:0]  img116;reg [7:0]  img117;reg [7:0]  img118;reg [7:0]  img119;reg [7:0]  img120;reg [7:0]  img121;reg [7:0]  img122;reg [7:0]  img123;reg [7:0]  img124;reg [7:0]  img125;reg [7:0]  img126;reg [7:0]  img127;reg [7:0]  img128;reg [7:0]  img129;reg [7:0]  img130;reg [7:0]  img131;reg [7:0]  img132;reg [7:0]  img133;reg [7:0]  img134;reg [7:0]  img135;reg [7:0]  img136;reg [7:0]  img137;reg [7:0]  img138;reg [7:0]  img139;reg [7:0]  img140;reg [7:0]  img141;reg [7:0]  img142;reg [7:0]  img143;reg [7:0]  img144;reg [7:0]  img145;reg [7:0]  img146;reg [7:0]  img147;reg [7:0]  img148;reg [7:0]  img149;reg [7:0]  img150;reg [7:0]  img151;reg [7:0]  img152;reg [7:0]  img153;reg [7:0]  img154;reg [7:0]  img155;reg [7:0]  img156;reg [7:0]  img157;reg [7:0]  img158;reg [7:0]  img159;reg [7:0]  img160;reg [7:0]  img161;reg [7:0]  img162;reg [7:0]  img163;reg [7:0]  img164;reg [7:0]  img165;reg [7:0]  img166;reg [7:0]  img167;reg [7:0]  img168;reg [7:0]  img169;reg [7:0]  img170;reg [7:0]  img171;reg [7:0]  img172;reg [7:0]  img173;reg [7:0]  img174;reg [7:0]  img175;reg [7:0]  img176;reg [7:0]  img177;reg [7:0]  img178;reg [7:0]  img179;reg [7:0]  img180;reg [7:0]  img181;reg [7:0]  img182;reg [7:0]  img183;reg [7:0]  img184;reg [7:0]  img185;reg [7:0]  img186;reg [7:0]  img187;reg [7:0]  img188;reg [7:0]  img189;reg [7:0]  img190;reg [7:0]  img191;reg [7:0]  img192;reg [7:0]  img193;reg [7:0]  img194;reg [7:0]  img195;reg [7:0]  img196;reg [7:0]  img197;reg [7:0]  img198;reg [7:0]  img199;reg [7:0]  img200;reg [7:0]  img201;reg [7:0]  img202;reg [7:0]  img203;reg [7:0]  img204;reg [7:0]  img205;reg [7:0]  img206;reg [7:0]  img207;reg [7:0]  img208;reg [7:0]  img209;reg [7:0]  img210;reg [7:0]  img211;reg [7:0]  img212;reg [7:0]  img213;reg [7:0]  img214;reg [7:0]  img215;reg [7:0]  img216;reg [7:0]  img217;reg [7:0]  img218;reg [7:0]  img219;reg [7:0]  img220;reg [7:0]  img221;reg [7:0]  img222;reg [7:0]  img223;reg [7:0]  img224;reg [7:0]  img225;reg [7:0]  img226;reg [7:0]  img227;reg [7:0]  img228;reg [7:0]  img229;reg [7:0]  img230;reg [7:0]  img231;reg [7:0]  img232;reg [7:0]  img233;reg [7:0]  img234;reg [7:0]  img235;reg [7:0]  img236;reg [7:0]  img237;reg [7:0]  img238;reg [7:0]  img239;reg [7:0]  img240;reg [7:0]  img241;reg [7:0]  img242;reg [7:0]  img243;reg [7:0]  img244;reg [7:0]  img245;reg [7:0]  img246;reg [7:0]  img247;reg [7:0]  img248;reg [7:0]  img249;reg [7:0]  img250;reg [7:0]  img251;reg [7:0]  img252;reg [7:0]  img253;reg [7:0]  img254;reg [7:0]  img255;reg [7:0]  img256;reg [7:0]  img257;reg [7:0]  img258;reg [7:0]  img259;reg [7:0]  img260;reg [7:0]  img261;reg [7:0]  img262;reg [7:0]  img263;reg [7:0]  img264;reg [7:0]  img265;reg [7:0]  img266;reg [7:0]  img267;reg [7:0]  img268;reg [7:0]  img269;reg [7:0]  img270;reg [7:0]  img271;reg [7:0]  img272;reg [7:0]  img273;reg [7:0]  img274;reg [7:0]  img275;reg [7:0]  img276;reg [7:0]  img277;reg [7:0]  img278;reg [7:0]  img279;reg [7:0]  img280;reg [7:0]  img281;reg [7:0]  img282;reg [7:0]  img283;reg [7:0]  img284;reg [7:0]  img285;reg [7:0]  img286;reg [7:0]  img287;reg [7:0]  img288;reg [7:0]  img289;reg [7:0]  img290;reg [7:0]  img291;reg [7:0]  img292;reg [7:0]  img293;reg [7:0]  img294;reg [7:0]  img295;reg [7:0]  img296;reg [7:0]  img297;reg [7:0]  img298;reg [7:0]  img299;reg [7:0]  img300;reg [7:0]  img301;reg [7:0]  img302;reg [7:0]  img303;reg [7:0]  img304;reg [7:0]  img305;reg [7:0]  img306;reg [7:0]  img307;reg [7:0]  img308;reg [7:0]  img309;reg [7:0]  img310;reg [7:0]  img311;reg [7:0]  img312;reg [7:0]  img313;reg [7:0]  img314;reg [7:0]  img315;reg [7:0]  img316;reg [7:0]  img317;reg [7:0]  img318;reg [7:0]  img319;reg [7:0]  img320;reg [7:0]  img321;reg [7:0]  img322;reg [7:0]  img323;reg [7:0]  img324;reg [7:0]  img325;reg [7:0]  img326;reg [7:0]  img327;reg [7:0]  img328;reg [7:0]  img329;reg [7:0]  img330;reg [7:0]  img331;reg [7:0]  img332;reg [7:0]  img333;reg [7:0]  img334;reg [7:0]  img335;reg [7:0]  img336;reg [7:0]  img337;reg [7:0]  img338;reg [7:0]  img339;reg [7:0]  img340;reg [7:0]  img341;reg [7:0]  img342;reg [7:0]  img343;reg [7:0]  img344;reg [7:0]  img345;reg [7:0]  img346;reg [7:0]  img347;reg [7:0]  img348;reg [7:0]  img349;reg [7:0]  img350;reg [7:0]  img351;reg [7:0]  img352;reg [7:0]  img353;reg [7:0]  img354;reg [7:0]  img355;reg [7:0]  img356;reg [7:0]  img357;reg [7:0]  img358;reg [7:0]  img359;reg [7:0]  img360;reg [7:0]  img361;reg [7:0]  img362;reg [7:0]  img363;reg [7:0]  img364;reg [7:0]  img365;reg [7:0]  img366;reg [7:0]  img367;reg [7:0]  img368;reg [7:0]  img369;reg [7:0]  img370;reg [7:0]  img371;reg [7:0]  img372;reg [7:0]  img373;reg [7:0]  img374;reg [7:0]  img375;reg [7:0]  img376;reg [7:0]  img377;reg [7:0]  img378;reg [7:0]  img379;reg [7:0]  img380;reg [7:0]  img381;reg [7:0]  img382;reg [7:0]  img383;reg [7:0]  img384;reg [7:0]  img385;reg [7:0]  img386;reg [7:0]  img387;reg [7:0]  img388;reg [7:0]  img389;reg [7:0]  img390;reg [7:0]  img391;reg [7:0]  img392;reg [7:0]  img393;reg [7:0]  img394;reg [7:0]  img395;reg [7:0]  img396;reg [7:0]  img397;reg [7:0]  img398;reg [7:0]  img399;reg [7:0]  img400;reg [7:0]  img401;reg [7:0]  img402;reg [7:0]  img403;reg [7:0]  img404;reg [7:0]  img405;reg [7:0]  img406;reg [7:0]  img407;reg [7:0]  img408;reg [7:0]  img409;reg [7:0]  img410;reg [7:0]  img411;reg [7:0]  img412;reg [7:0]  img413;reg [7:0]  img414;reg [7:0]  img415;reg [7:0]  img416;reg [7:0]  img417;reg [7:0]  img418;reg [7:0]  img419;reg [7:0]  img420;reg [7:0]  img421;reg [7:0]  img422;reg [7:0]  img423;reg [7:0]  img424;reg [7:0]  img425;reg [7:0]  img426;reg [7:0]  img427;reg [7:0]  img428;reg [7:0]  img429;reg [7:0]  img430;reg [7:0]  img431;reg [7:0]  img432;reg [7:0]  img433;reg [7:0]  img434;reg [7:0]  img435;reg [7:0]  img436;reg [7:0]  img437;reg [7:0]  img438;reg [7:0]  img439;reg [7:0]  img440;reg [7:0]  img441;reg [7:0]  img442;reg [7:0]  img443;reg [7:0]  img444;reg [7:0]  img445;reg [7:0]  img446;reg [7:0]  img447;reg [7:0]  img448;reg [7:0]  img449;reg [7:0]  img450;reg [7:0]  img451;reg [7:0]  img452;reg [7:0]  img453;reg [7:0]  img454;reg [7:0]  img455;reg [7:0]  img456;reg [7:0]  img457;reg [7:0]  img458;reg [7:0]  img459;reg [7:0]  img460;reg [7:0]  img461;reg [7:0]  img462;reg [7:0]  img463;reg [7:0]  img464;reg [7:0]  img465;reg [7:0]  img466;reg [7:0]  img467;reg [7:0]  img468;reg [7:0]  img469;reg [7:0]  img470;reg [7:0]  img471;reg [7:0]  img472;reg [7:0]  img473;reg [7:0]  img474;reg [7:0]  img475;reg [7:0]  img476;reg [7:0]  img477;reg [7:0]  img478;reg [7:0]  img479;reg [7:0]  img480;reg [7:0]  img481;reg [7:0]  img482;reg [7:0]  img483;reg [7:0]  img484;reg [7:0]  img485;reg [7:0]  img486;reg [7:0]  img487;reg [7:0]  img488;reg [7:0]  img489;reg [7:0]  img490;reg [7:0]  img491;reg [7:0]  img492;reg [7:0]  img493;reg [7:0]  img494;reg [7:0]  img495;reg [7:0]  img496;reg [7:0]  img497;reg [7:0]  img498;reg [7:0]  img499;reg [7:0]  img500;reg [7:0]  img501;reg [7:0]  img502;reg [7:0]  img503;reg [7:0]  img504;reg [7:0]  img505;reg [7:0]  img506;reg [7:0]  img507;reg [7:0]  img508;reg [7:0]  img509;reg [7:0]  img510;reg [7:0]  img511;reg [7:0]  img512;reg [7:0]  img513;reg [7:0]  img514;reg [7:0]  img515;reg [7:0]  img516;reg [7:0]  img517;reg [7:0]  img518;reg [7:0]  img519;reg [7:0]  img520;reg [7:0]  img521;reg [7:0]  img522;reg [7:0]  img523;reg [7:0]  img524;reg [7:0]  img525;reg [7:0]  img526;reg [7:0]  img527;reg [7:0]  img528;reg [7:0]  img529;reg [7:0]  img530;reg [7:0]  img531;reg [7:0]  img532;reg [7:0]  img533;reg [7:0]  img534;reg [7:0]  img535;reg [7:0]  img536;reg [7:0]  img537;reg [7:0]  img538;reg [7:0]  img539;reg [7:0]  img540;reg [7:0]  img541;reg [7:0]  img542;reg [7:0]  img543;reg [7:0]  img544;reg [7:0]  img545;reg [7:0]  img546;reg [7:0]  img547;reg [7:0]  img548;reg [7:0]  img549;reg [7:0]  img550;reg [7:0]  img551;reg [7:0]  img552;reg [7:0]  img553;reg [7:0]  img554;reg [7:0]  img555;reg [7:0]  img556;reg [7:0]  img557;reg [7:0]  img558;reg [7:0]  img559;reg [7:0]  img560;reg [7:0]  img561;reg [7:0]  img562;reg [7:0]  img563;reg [7:0]  img564;reg [7:0]  img565;reg [7:0]  img566;reg [7:0]  img567;reg [7:0]  img568;reg [7:0]  img569;reg [7:0]  img570;reg [7:0]  img571;reg [7:0]  img572;reg [7:0]  img573;reg [7:0]  img574;reg [7:0]  img575;reg [7:0]  img576;reg [7:0]  img577;reg [7:0]  img578;reg [7:0]  img579;reg [7:0]  img580;reg [7:0]  img581;reg [7:0]  img582;reg [7:0]  img583;reg [7:0]  img584;reg [7:0]  img585;reg [7:0]  img586;reg [7:0]  img587;reg [7:0]  img588;reg [7:0]  img589;reg [7:0]  img590;reg [7:0]  img591;reg [7:0]  img592;reg [7:0]  img593;reg [7:0]  img594;reg [7:0]  img595;reg [7:0]  img596;reg [7:0]  img597;reg [7:0]  img598;reg [7:0]  img599;reg [7:0]  img600;reg [7:0]  img601;reg [7:0]  img602;reg [7:0]  img603;reg [7:0]  img604;reg [7:0]  img605;reg [7:0]  img606;reg [7:0]  img607;reg [7:0]  img608;reg [7:0]  img609;reg [7:0]  img610;reg [7:0]  img611;reg [7:0]  img612;reg [7:0]  img613;reg [7:0]  img614;reg [7:0]  img615;reg [7:0]  img616;reg [7:0]  img617;reg [7:0]  img618;reg [7:0]  img619;reg [7:0]  img620;reg [7:0]  img621;reg [7:0]  img622;reg [7:0]  img623;reg [7:0]  img624;reg [7:0]  img625;reg [7:0]  img626;reg [7:0]  img627;reg [7:0]  img628;reg [7:0]  img629;reg [7:0]  img630;reg [7:0]  img631;reg [7:0]  img632;reg [7:0]  img633;reg [7:0]  img634;reg [7:0]  img635;reg [7:0]  img636;reg [7:0]  img637;reg [7:0]  img638;reg [7:0]  img639;reg [7:0]  img640;reg [7:0]  img641;reg [7:0]  img642;reg [7:0]  img643;reg [7:0]  img644;reg [7:0]  img645;reg [7:0]  img646;reg [7:0]  img647;reg [7:0]  img648;reg [7:0]  img649;reg [7:0]  img650;reg [7:0]  img651;reg [7:0]  img652;reg [7:0]  img653;reg [7:0]  img654;reg [7:0]  img655;reg [7:0]  img656;reg [7:0]  img657;reg [7:0]  img658;reg [7:0]  img659;reg [7:0]  img660;reg [7:0]  img661;reg [7:0]  img662;reg [7:0]  img663;reg [7:0]  img664;reg [7:0]  img665;reg [7:0]  img666;reg [7:0]  img667;reg [7:0]  img668;reg [7:0]  img669;reg [7:0]  img670;reg [7:0]  img671;reg [7:0]  img672;reg [7:0]  img673;reg [7:0]  img674;reg [7:0]  img675;reg [7:0]  img676;reg [7:0]  img677;reg [7:0]  img678;reg [7:0]  img679;reg [7:0]  img680;reg [7:0]  img681;reg [7:0]  img682;reg [7:0]  img683;reg [7:0]  img684;reg [7:0]  img685;reg [7:0]  img686;reg [7:0]  img687;reg [7:0]  img688;reg [7:0]  img689;reg [7:0]  img690;reg [7:0]  img691;reg [7:0]  img692;reg [7:0]  img693;reg [7:0]  img694;reg [7:0]  img695;reg [7:0]  img696;reg [7:0]  img697;reg [7:0]  img698;reg [7:0]  img699;reg [7:0]  img700;reg [7:0]  img701;reg [7:0]  img702;reg [7:0]  img703;reg [7:0]  img704;reg [7:0]  img705;reg [7:0]  img706;reg [7:0]  img707;reg [7:0]  img708;reg [7:0]  img709;reg [7:0]  img710;reg [7:0]  img711;reg [7:0]  img712;reg [7:0]  img713;reg [7:0]  img714;reg [7:0]  img715;reg [7:0]  img716;reg [7:0]  img717;reg [7:0]  img718;reg [7:0]  img719;reg [7:0]  img720;reg [7:0]  img721;reg [7:0]  img722;reg [7:0]  img723;reg [7:0]  img724;reg [7:0]  img725;reg [7:0]  img726;reg [7:0]  img727;reg [7:0]  img728;reg [7:0]  img729;reg [7:0]  img730;reg [7:0]  img731;reg [7:0]  img732;reg [7:0]  img733;reg [7:0]  img734;reg [7:0]  img735;reg [7:0]  img736;reg [7:0]  img737;reg [7:0]  img738;reg [7:0]  img739;reg [7:0]  img740;reg [7:0]  img741;reg [7:0]  img742;reg [7:0]  img743;reg [7:0]  img744;reg [7:0]  img745;reg [7:0]  img746;reg [7:0]  img747;reg [7:0]  img748;reg [7:0]  img749;reg [7:0]  img750;reg [7:0]  img751;reg [7:0]  img752;reg [7:0]  img753;reg [7:0]  img754;reg [7:0]  img755;reg [7:0]  img756;reg [7:0]  img757;reg [7:0]  img758;reg [7:0]  img759;reg [7:0]  img760;reg [7:0]  img761;reg [7:0]  img762;reg [7:0]  img763;reg [7:0]  img764;reg [7:0]  img765;reg [7:0]  img766;reg [7:0]  img767;reg [7:0]  img768;reg [7:0]  img769;reg [7:0]  img770;reg [7:0]  img771;reg [7:0]  img772;reg [7:0]  img773;reg [7:0]  img774;reg [7:0]  img775;reg [7:0]  img776;reg [7:0]  img777;reg [7:0]  img778;reg [7:0]  img779;reg [7:0]  img780;reg [7:0]  img781;reg [7:0]  img782;reg [7:0]  img783;
wire [3:0] predict;
       net #(64,2,784) 
       UDT
      (.clk(clk),
       .rst(rst),
        .img0(img0),.img1(img1),.img2(img2),.img3(img3),.img4(img4),.img5(img5),.img6(img6),.img7(img7),.img8(img8),.img9(img9),.img10(img10),.img11(img11),.img12(img12),.img13(img13),.img14(img14),.img15(img15),.img16(img16),.img17(img17),.img18(img18),.img19(img19),.img20(img20),.img21(img21),.img22(img22),.img23(img23),.img24(img24),.img25(img25),.img26(img26),.img27(img27),.img28(img28),.img29(img29),.img30(img30),.img31(img31),.img32(img32),.img33(img33),.img34(img34),.img35(img35),.img36(img36),.img37(img37),.img38(img38),.img39(img39),.img40(img40),.img41(img41),.img42(img42),.img43(img43),.img44(img44),.img45(img45),.img46(img46),.img47(img47),.img48(img48),.img49(img49),.img50(img50),.img51(img51),.img52(img52),.img53(img53),.img54(img54),.img55(img55),.img56(img56),.img57(img57),.img58(img58),.img59(img59),.img60(img60),.img61(img61),.img62(img62),.img63(img63),.img64(img64),.img65(img65),.img66(img66),.img67(img67),.img68(img68),.img69(img69),.img70(img70),.img71(img71),.img72(img72),.img73(img73),.img74(img74),.img75(img75),.img76(img76),.img77(img77),.img78(img78),.img79(img79),.img80(img80),.img81(img81),.img82(img82),.img83(img83),.img84(img84),.img85(img85),.img86(img86),.img87(img87),.img88(img88),.img89(img89),.img90(img90),.img91(img91),.img92(img92),.img93(img93),.img94(img94),.img95(img95),.img96(img96),.img97(img97),.img98(img98),.img99(img99),.img100(img100),.img101(img101),.img102(img102),.img103(img103),.img104(img104),.img105(img105),.img106(img106),.img107(img107),.img108(img108),.img109(img109),.img110(img110),.img111(img111),.img112(img112),.img113(img113),.img114(img114),.img115(img115),.img116(img116),.img117(img117),.img118(img118),.img119(img119),.img120(img120),.img121(img121),.img122(img122),.img123(img123),.img124(img124),.img125(img125),.img126(img126),.img127(img127),.img128(img128),.img129(img129),.img130(img130),.img131(img131),.img132(img132),.img133(img133),.img134(img134),.img135(img135),.img136(img136),.img137(img137),.img138(img138),.img139(img139),.img140(img140),.img141(img141),.img142(img142),.img143(img143),.img144(img144),.img145(img145),.img146(img146),.img147(img147),.img148(img148),.img149(img149),.img150(img150),.img151(img151),.img152(img152),.img153(img153),.img154(img154),.img155(img155),.img156(img156),.img157(img157),.img158(img158),.img159(img159),.img160(img160),.img161(img161),.img162(img162),.img163(img163),.img164(img164),.img165(img165),.img166(img166),.img167(img167),.img168(img168),.img169(img169),.img170(img170),.img171(img171),.img172(img172),.img173(img173),.img174(img174),.img175(img175),.img176(img176),.img177(img177),.img178(img178),.img179(img179),.img180(img180),.img181(img181),.img182(img182),.img183(img183),.img184(img184),.img185(img185),.img186(img186),.img187(img187),.img188(img188),.img189(img189),.img190(img190),.img191(img191),.img192(img192),.img193(img193),.img194(img194),.img195(img195),.img196(img196),.img197(img197),.img198(img198),.img199(img199),.img200(img200),.img201(img201),.img202(img202),.img203(img203),.img204(img204),.img205(img205),.img206(img206),.img207(img207),.img208(img208),.img209(img209),.img210(img210),.img211(img211),.img212(img212),.img213(img213),.img214(img214),.img215(img215),.img216(img216),.img217(img217),.img218(img218),.img219(img219),.img220(img220),.img221(img221),.img222(img222),.img223(img223),.img224(img224),.img225(img225),.img226(img226),.img227(img227),.img228(img228),.img229(img229),.img230(img230),.img231(img231),.img232(img232),.img233(img233),.img234(img234),.img235(img235),.img236(img236),.img237(img237),.img238(img238),.img239(img239),.img240(img240),.img241(img241),.img242(img242),.img243(img243),.img244(img244),.img245(img245),.img246(img246),.img247(img247),.img248(img248),.img249(img249),.img250(img250),.img251(img251),.img252(img252),.img253(img253),.img254(img254),.img255(img255),.img256(img256),.img257(img257),.img258(img258),.img259(img259),.img260(img260),.img261(img261),.img262(img262),.img263(img263),.img264(img264),.img265(img265),.img266(img266),.img267(img267),.img268(img268),.img269(img269),.img270(img270),.img271(img271),.img272(img272),.img273(img273),.img274(img274),.img275(img275),.img276(img276),.img277(img277),.img278(img278),.img279(img279),.img280(img280),.img281(img281),.img282(img282),.img283(img283),.img284(img284),.img285(img285),.img286(img286),.img287(img287),.img288(img288),.img289(img289),.img290(img290),.img291(img291),.img292(img292),.img293(img293),.img294(img294),.img295(img295),.img296(img296),.img297(img297),.img298(img298),.img299(img299),.img300(img300),.img301(img301),.img302(img302),.img303(img303),.img304(img304),.img305(img305),.img306(img306),.img307(img307),.img308(img308),.img309(img309),.img310(img310),.img311(img311),.img312(img312),.img313(img313),.img314(img314),.img315(img315),.img316(img316),.img317(img317),.img318(img318),.img319(img319),.img320(img320),.img321(img321),.img322(img322),.img323(img323),.img324(img324),.img325(img325),.img326(img326),.img327(img327),.img328(img328),.img329(img329),.img330(img330),.img331(img331),.img332(img332),.img333(img333),.img334(img334),.img335(img335),.img336(img336),.img337(img337),.img338(img338),.img339(img339),.img340(img340),.img341(img341),.img342(img342),.img343(img343),.img344(img344),.img345(img345),.img346(img346),.img347(img347),.img348(img348),.img349(img349),.img350(img350),.img351(img351),.img352(img352),.img353(img353),.img354(img354),.img355(img355),.img356(img356),.img357(img357),.img358(img358),.img359(img359),.img360(img360),.img361(img361),.img362(img362),.img363(img363),.img364(img364),.img365(img365),.img366(img366),.img367(img367),.img368(img368),.img369(img369),.img370(img370),.img371(img371),.img372(img372),.img373(img373),.img374(img374),.img375(img375),.img376(img376),.img377(img377),.img378(img378),.img379(img379),.img380(img380),.img381(img381),.img382(img382),.img383(img383),.img384(img384),.img385(img385),.img386(img386),.img387(img387),.img388(img388),.img389(img389),.img390(img390),.img391(img391),.img392(img392),.img393(img393),.img394(img394),.img395(img395),.img396(img396),.img397(img397),.img398(img398),.img399(img399),.img400(img400),.img401(img401),.img402(img402),.img403(img403),.img404(img404),.img405(img405),.img406(img406),.img407(img407),.img408(img408),.img409(img409),.img410(img410),.img411(img411),.img412(img412),.img413(img413),.img414(img414),.img415(img415),.img416(img416),.img417(img417),.img418(img418),.img419(img419),.img420(img420),.img421(img421),.img422(img422),.img423(img423),.img424(img424),.img425(img425),.img426(img426),.img427(img427),.img428(img428),.img429(img429),.img430(img430),.img431(img431),.img432(img432),.img433(img433),.img434(img434),.img435(img435),.img436(img436),.img437(img437),.img438(img438),.img439(img439),.img440(img440),.img441(img441),.img442(img442),.img443(img443),.img444(img444),.img445(img445),.img446(img446),.img447(img447),.img448(img448),.img449(img449),.img450(img450),.img451(img451),.img452(img452),.img453(img453),.img454(img454),.img455(img455),.img456(img456),.img457(img457),.img458(img458),.img459(img459),.img460(img460),.img461(img461),.img462(img462),.img463(img463),.img464(img464),.img465(img465),.img466(img466),.img467(img467),.img468(img468),.img469(img469),.img470(img470),.img471(img471),.img472(img472),.img473(img473),.img474(img474),.img475(img475),.img476(img476),.img477(img477),.img478(img478),.img479(img479),.img480(img480),.img481(img481),.img482(img482),.img483(img483),.img484(img484),.img485(img485),.img486(img486),.img487(img487),.img488(img488),.img489(img489),.img490(img490),.img491(img491),.img492(img492),.img493(img493),.img494(img494),.img495(img495),.img496(img496),.img497(img497),.img498(img498),.img499(img499),.img500(img500),.img501(img501),.img502(img502),.img503(img503),.img504(img504),.img505(img505),.img506(img506),.img507(img507),.img508(img508),.img509(img509),.img510(img510),.img511(img511),.img512(img512),.img513(img513),.img514(img514),.img515(img515),.img516(img516),.img517(img517),.img518(img518),.img519(img519),.img520(img520),.img521(img521),.img522(img522),.img523(img523),.img524(img524),.img525(img525),.img526(img526),.img527(img527),.img528(img528),.img529(img529),.img530(img530),.img531(img531),.img532(img532),.img533(img533),.img534(img534),.img535(img535),.img536(img536),.img537(img537),.img538(img538),.img539(img539),.img540(img540),.img541(img541),.img542(img542),.img543(img543),.img544(img544),.img545(img545),.img546(img546),.img547(img547),.img548(img548),.img549(img549),.img550(img550),.img551(img551),.img552(img552),.img553(img553),.img554(img554),.img555(img555),.img556(img556),.img557(img557),.img558(img558),.img559(img559),.img560(img560),.img561(img561),.img562(img562),.img563(img563),.img564(img564),.img565(img565),.img566(img566),.img567(img567),.img568(img568),.img569(img569),.img570(img570),.img571(img571),.img572(img572),.img573(img573),.img574(img574),.img575(img575),.img576(img576),.img577(img577),.img578(img578),.img579(img579),.img580(img580),.img581(img581),.img582(img582),.img583(img583),.img584(img584),.img585(img585),.img586(img586),.img587(img587),.img588(img588),.img589(img589),.img590(img590),.img591(img591),.img592(img592),.img593(img593),.img594(img594),.img595(img595),.img596(img596),.img597(img597),.img598(img598),.img599(img599),.img600(img600),.img601(img601),.img602(img602),.img603(img603),.img604(img604),.img605(img605),.img606(img606),.img607(img607),.img608(img608),.img609(img609),.img610(img610),.img611(img611),.img612(img612),.img613(img613),.img614(img614),.img615(img615),.img616(img616),.img617(img617),.img618(img618),.img619(img619),.img620(img620),.img621(img621),.img622(img622),.img623(img623),.img624(img624),.img625(img625),.img626(img626),.img627(img627),.img628(img628),.img629(img629),.img630(img630),.img631(img631),.img632(img632),.img633(img633),.img634(img634),.img635(img635),.img636(img636),.img637(img637),.img638(img638),.img639(img639),.img640(img640),.img641(img641),.img642(img642),.img643(img643),.img644(img644),.img645(img645),.img646(img646),.img647(img647),.img648(img648),.img649(img649),.img650(img650),.img651(img651),.img652(img652),.img653(img653),.img654(img654),.img655(img655),.img656(img656),.img657(img657),.img658(img658),.img659(img659),.img660(img660),.img661(img661),.img662(img662),.img663(img663),.img664(img664),.img665(img665),.img666(img666),.img667(img667),.img668(img668),.img669(img669),.img670(img670),.img671(img671),.img672(img672),.img673(img673),.img674(img674),.img675(img675),.img676(img676),.img677(img677),.img678(img678),.img679(img679),.img680(img680),.img681(img681),.img682(img682),.img683(img683),.img684(img684),.img685(img685),.img686(img686),.img687(img687),.img688(img688),.img689(img689),.img690(img690),.img691(img691),.img692(img692),.img693(img693),.img694(img694),.img695(img695),.img696(img696),.img697(img697),.img698(img698),.img699(img699),.img700(img700),.img701(img701),.img702(img702),.img703(img703),.img704(img704),.img705(img705),.img706(img706),.img707(img707),.img708(img708),.img709(img709),.img710(img710),.img711(img711),.img712(img712),.img713(img713),.img714(img714),.img715(img715),.img716(img716),.img717(img717),.img718(img718),.img719(img719),.img720(img720),.img721(img721),.img722(img722),.img723(img723),.img724(img724),.img725(img725),.img726(img726),.img727(img727),.img728(img728),.img729(img729),.img730(img730),.img731(img731),.img732(img732),.img733(img733),.img734(img734),.img735(img735),.img736(img736),.img737(img737),.img738(img738),.img739(img739),.img740(img740),.img741(img741),.img742(img742),.img743(img743),.img744(img744),.img745(img745),.img746(img746),.img747(img747),.img748(img748),.img749(img749),.img750(img750),.img751(img751),.img752(img752),.img753(img753),.img754(img754),.img755(img755),.img756(img756),.img757(img757),.img758(img758),.img759(img759),.img760(img760),.img761(img761),.img762(img762),.img763(img763),.img764(img764),.img765(img765),.img766(img766),.img767(img767),.img768(img768),.img769(img769),.img770(img770),.img771(img771),.img772(img772),.img773(img773),.img774(img774),.img775(img775),.img776(img776),.img777(img777),.img778(img778),.img779(img779),.img780(img780),.img781(img781),.img782(img782),.img783(img783),
       .predict(predict)
       );
always #5 clk=~clk;
reg[3:0] read_data [0:100];
integer i,hit;

initial 
   begin
       i=-4;hit=0;
       $display("begin read label file... ");
       $readmemh("label.mem",read_data);
   end
always@(posedge clk)
   begin
       $display("data     :%d predict    :%d",read_data[i],predict); 
           if(predict==read_data[i])
               begin
                   hit=hit+1;
               end
       i=i+1'b1;
   end
initial 
begin
rst=1'b1;clk=1'b0;

#10 rst=1'b0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd42;img203=8'd93;img204=8'd80;img205=8'd76;img206=8'd30;img207=8'd18;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd111;img231=8'd127;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd121;img236=8'd99;img237=8'd99;img238=8'd99;img239=8'd99;img240=8'd99;img241=8'd99;img242=8'd99;img243=8'd99;img244=8'd85;img245=8'd26;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd34;img259=8'd57;img260=8'd36;img261=8'd57;img262=8'd82;img263=8'd114;img264=8'd127;img265=8'd113;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd125;img270=8'd115;img271=8'd127;img272=8'd127;img273=8'd70;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd9;img292=8'd33;img293=8'd7;img294=8'd34;img295=8'd34;img296=8'd34;img297=8'd30;img298=8'd11;img299=8'd118;img300=8'd127;img301=8'd53;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd42;img327=8'd127;img328=8'd105;img329=8'd9;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd11;img354=8'd117;img355=8'd128;img356=8'd42;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd65;img382=8'd127;img383=8'd119;img384=8'd22;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd30;img409=8'd125;img410=8'd127;img411=8'd31;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd67;img437=8'd127;img438=8'd94;img439=8'd3;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd5;img464=8'd103;img465=8'd124;img466=8'd29;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd63;img492=8'd127;img493=8'd91;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd38;img519=8'd126;img520=8'd120;img521=8'd29;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd10;img546=8'd111;img547=8'd127;img548=8'd83;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd2;img573=8'd102;img574=8'd127;img575=8'd110;img576=8'd18;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd19;img601=8'd127;img602=8'd127;img603=8'd39;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd16;img628=8'd112;img629=8'd127;img630=8'd58;img631=8'd1;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd67;img656=8'd127;img657=8'd127;img658=8'd26;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd31;img683=8'd121;img684=8'd127;img685=8'd127;img686=8'd26;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd61;img711=8'd127;img712=8'd127;img713=8'd110;img714=8'd20;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd61;img739=8'd127;img740=8'd104;img741=8'd9;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd58;img95=8'd63;img96=8'd86;img97=8'd128;img98=8'd128;img99=8'd75;img100=8'd47;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd85;img122=8'd127;img123=8'd127;img124=8'd127;img125=8'd127;img126=8'd127;img127=8'd127;img128=8'd109;img129=8'd15;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd85;img149=8'd127;img150=8'd127;img151=8'd127;img152=8'd107;img153=8'd71;img154=8'd88;img155=8'd127;img156=8'd127;img157=8'd61;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd26;img176=8'd125;img177=8'd127;img178=8'd105;img179=8'd16;img180=8'd6;img181=8'd0;img182=8'd3;img183=8'd103;img184=8'd127;img185=8'd70;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd39;img204=8'd126;img205=8'd105;img206=8'd13;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd61;img211=8'd124;img212=8'd127;img213=8'd33;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd16;img233=8'd9;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd105;img239=8'd127;img240=8'd127;img241=8'd33;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd59;img266=8'd124;img267=8'd127;img268=8'd99;img269=8'd5;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd38;img293=8'd124;img294=8'd127;img295=8'd116;img296=8'd32;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd64;img321=8'd127;img322=8'd127;img323=8'd72;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd88;img348=8'd123;img349=8'd127;img350=8'd80;img351=8'd6;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd13;img375=8'd117;img376=8'd127;img377=8'd117;img378=8'd18;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd99;img403=8'd127;img404=8'd127;img405=8'd71;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd39;img430=8'd124;img431=8'd127;img432=8'd95;img433=8'd6;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd10;img457=8'd100;img458=8'd127;img459=8'd127;img460=8'd71;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd67;img485=8'd127;img486=8'd127;img487=8'd87;img488=8'd6;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd124;img513=8'd127;img514=8'd127;img515=8'd13;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd124;img541=8'd127;img542=8'd127;img543=8'd22;img544=8'd10;img545=8'd10;img546=8'd10;img547=8'd10;img548=8'd3;img549=8'd0;img550=8'd3;img551=8'd10;img552=8'd10;img553=8'd19;img554=8'd75;img555=8'd75;img556=8'd75;img557=8'd74;img558=8'd5;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd124;img569=8'd127;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd84;img577=8'd72;img578=8'd83;img579=8'd127;img580=8'd127;img581=8'd127;img582=8'd127;img583=8'd127;img584=8'd127;img585=8'd127;img586=8'd62;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd87;img597=8'd127;img598=8'd127;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd127;img607=8'd127;img608=8'd125;img609=8'd124;img610=8'd124;img611=8'd85;img612=8'd59;img613=8'd59;img614=8'd29;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd59;img626=8'd62;img627=8'd62;img628=8'd62;img629=8'd83;img630=8'd127;img631=8'd127;img632=8'd127;img633=8'd78;img634=8'd62;img635=8'd62;img636=8'd21;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd19;img129=8'd127;img130=8'd55;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd44;img157=8'd126;img158=8'd41;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd68;img185=8'd121;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd23;img212=8'd122;img213=8'd75;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd42;img240=8'd127;img241=8'd32;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd101;img268=8'd112;img269=8'd6;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd16;img295=8'd127;img296=8'd108;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd48;img323=8'd127;img324=8'd98;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd70;img351=8'd127;img352=8'd39;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd29;img378=8'd119;img379=8'd103;img380=8'd4;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd62;img406=8'd128;img407=8'd83;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd86;img434=8'd127;img435=8'd41;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd12;img461=8'd116;img462=8'd108;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd60;img489=8'd127;img490=8'd80;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd76;img517=8'd127;img518=8'd71;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd114;img545=8'd127;img546=8'd33;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd31;img572=8'd126;img573=8'd127;img574=8'd33;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd71;img600=8'd127;img601=8'd103;img602=8'd2;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd5;img627=8'd108;img628=8'd127;img629=8'd61;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd3;img655=8'd99;img656=8'd88;img657=8'd5;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd6;img125=8'd75;img126=8'd127;img127=8'd101;img128=8'd16;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd19;img153=8'd126;img154=8'd126;img155=8'd127;img156=8'd54;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd11;img180=8'd99;img181=8'd126;img182=8'd126;img183=8'd127;img184=8'd54;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd55;img207=8'd95;img208=8'd126;img209=8'd126;img210=8'd126;img211=8'd127;img212=8'd85;img213=8'd55;img214=8'd31;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd127;img235=8'd126;img236=8'd126;img237=8'd126;img238=8'd126;img239=8'd127;img240=8'd126;img241=8'd126;img242=8'd110;img243=8'd26;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd91;img262=8'd128;img263=8'd127;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd117;img268=8'd111;img269=8'd127;img270=8'd127;img271=8'd127;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd32;img289=8'd111;img290=8'd127;img291=8'd126;img292=8'd126;img293=8'd126;img294=8'd74;img295=8'd39;img296=8'd31;img297=8'd64;img298=8'd126;img299=8'd126;img300=8'd53;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd16;img316=8'd116;img317=8'd126;img318=8'd127;img319=8'd126;img320=8'd110;img321=8'd69;img322=8'd5;img323=8'd0;img324=8'd0;img325=8'd16;img326=8'd115;img327=8'd126;img328=8'd122;img329=8'd57;img330=8'd3;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd19;img344=8'd126;img345=8'd126;img346=8'd127;img347=8'd94;img348=8'd10;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd55;img355=8'd126;img356=8'd127;img357=8'd126;img358=8'd18;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd19;img372=8'd126;img373=8'd126;img374=8'd101;img375=8'd15;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd16;img383=8'd100;img384=8'd127;img385=8'd126;img386=8'd18;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd19;img400=8'd127;img401=8'd127;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd16;img411=8'd101;img412=8'd128;img413=8'd127;img414=8'd82;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd70;img428=8'd126;img429=8'd126;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd55;img439=8'd126;img440=8'd127;img441=8'd126;img442=8'd18;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd109;img456=8'd126;img457=8'd126;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd11;img465=8'd32;img466=8'd116;img467=8'd126;img468=8'd127;img469=8'd115;img470=8'd15;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd109;img484=8'd126;img485=8'd126;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd72;img493=8'd126;img494=8'd126;img495=8'd126;img496=8'd111;img497=8'd31;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd109;img512=8'd126;img513=8'd126;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd91;img520=8'd111;img521=8'd126;img522=8'd126;img523=8'd126;img524=8'd90;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd109;img540=8'd127;img541=8'd127;img542=8'd37;img543=8'd37;img544=8'd114;img545=8'd127;img546=8'd127;img547=8'd128;img548=8'd127;img549=8'd127;img550=8'd127;img551=8'd127;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd57;img568=8'd126;img569=8'd126;img570=8'd127;img571=8'd126;img572=8'd126;img573=8'd126;img574=8'd126;img575=8'd127;img576=8'd126;img577=8'd126;img578=8'd126;img579=8'd74;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd16;img596=8'd115;img597=8'd126;img598=8'd127;img599=8'd126;img600=8'd126;img601=8'd126;img602=8'd126;img603=8'd127;img604=8'd115;img605=8'd95;img606=8'd18;img607=8'd5;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd31;img625=8'd71;img626=8'd127;img627=8'd126;img628=8'd126;img629=8'd126;img630=8'd126;img631=8'd127;img632=8'd54;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd36;img655=8'd87;img656=8'd126;img657=8'd87;img658=8'd36;img659=8'd36;img660=8'd15;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd25;img151=8'd112;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd35;img160=8'd15;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd61;img179=8'd116;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd74;img188=8'd84;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd2;img206=8'd98;img207=8'd116;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd48;img216=8'd105;img217=8'd6;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd35;img234=8'd126;img235=8'd67;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd57;img244=8'd126;img245=8'd11;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd23;img261=8'd118;img262=8'd109;img263=8'd6;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd96;img272=8'd126;img273=8'd11;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd84;img289=8'd124;img290=8'd27;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd9;img299=8'd128;img300=8'd127;img301=8'd11;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd42;img316=8'd121;img317=8'd106;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd71;img327=8'd127;img328=8'd95;img329=8'd3;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd85;img344=8'd126;img345=8'd53;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd16;img354=8'd116;img355=8'd125;img356=8'd33;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd8;img371=8'd113;img372=8'd126;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd67;img382=8'd126;img383=8'd106;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd11;img399=8'd126;img400=8'd82;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd85;img410=8'd126;img411=8'd84;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd5;img427=8'd102;img428=8'd105;img429=8'd9;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd11;img437=8'd127;img438=8'd127;img439=8'd54;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd85;img456=8'd126;img457=8'd100;img458=8'd43;img459=8'd43;img460=8'd43;img461=8'd43;img462=8'd65;img463=8'd82;img464=8'd98;img465=8'd126;img466=8'd126;img467=8'd53;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd21;img484=8'd85;img485=8'd123;img486=8'd126;img487=8'd126;img488=8'd126;img489=8'd126;img490=8'd116;img491=8'd116;img492=8'd126;img493=8'd126;img494=8'd126;img495=8'd5;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd25;img514=8'd42;img515=8'd42;img516=8'd42;img517=8'd42;img518=8'd0;img519=8'd0;img520=8'd81;img521=8'd126;img522=8'd126;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd64;img549=8'd126;img550=8'd126;img551=8'd23;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd64;img577=8'd127;img578=8'd127;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd64;img605=8'd126;img606=8'd126;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd68;img633=8'd126;img634=8'd122;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd116;img661=8'd118;img662=8'd56;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd90;img689=8'd33;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd39;img157=8'd127;img158=8'd54;img159=8'd2;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd10;img184=8'd114;img185=8'd127;img186=8'd127;img187=8'd5;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd41;img212=8'd127;img213=8'd127;img214=8'd83;img215=8'd1;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd4;img239=8'd102;img240=8'd127;img241=8'd127;img242=8'd37;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd27;img267=8'd127;img268=8'd127;img269=8'd125;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd67;img295=8'd127;img296=8'd127;img297=8'd90;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd98;img323=8'd127;img324=8'd124;img325=8'd24;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd29;img350=8'd127;img351=8'd127;img352=8'd119;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd56;img378=8'd127;img379=8'd127;img380=8'd66;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd82;img406=8'd127;img407=8'd119;img408=8'd14;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd30;img433=8'd126;img434=8'd127;img435=8'd112;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd40;img461=8'd127;img462=8'd127;img463=8'd77;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd82;img489=8'd127;img490=8'd119;img491=8'd27;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd14;img516=8'd126;img517=8'd127;img518=8'd105;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd43;img544=8'd127;img545=8'd127;img546=8'd66;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd53;img572=8'd127;img573=8'd117;img574=8'd10;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd88;img600=8'd127;img601=8'd102;img602=8'd3;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd3;img627=8'd106;img628=8'd127;img629=8'd98;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd2;img655=8'd79;img656=8'd127;img657=8'd80;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd13;img684=8'd79;img685=8'd54;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd11;img150=8'd96;img151=8'd67;img152=8'd16;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd8;img162=8'd39;img163=8'd3;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd9;img177=8'd118;img178=8'd125;img179=8'd85;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd8;img189=8'd110;img190=8'd121;img191=8'd19;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd10;img204=8'd95;img205=8'd127;img206=8'd74;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd70;img217=8'd127;img218=8'd50;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd35;img232=8'd127;img233=8'd127;img234=8'd11;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd22;img244=8'd127;img245=8'd87;img246=8'd7;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd11;img259=8'd77;img260=8'd127;img261=8'd48;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd22;img271=8'd116;img272=8'd127;img273=8'd46;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd82;img287=8'd128;img288=8'd102;img289=8'd6;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd52;img299=8'd127;img300=8'd79;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd81;img315=8'd127;img316=8'd89;img317=8'd3;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd5;img325=8'd66;img326=8'd119;img327=8'd127;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd81;img343=8'd127;img344=8'd127;img345=8'd96;img346=8'd88;img347=8'd35;img348=8'd35;img349=8'd35;img350=8'd35;img351=8'd67;img352=8'd99;img353=8'd127;img354=8'd127;img355=8'd85;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd26;img371=8'd114;img372=8'd127;img373=8'd127;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd110;img383=8'd18;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd9;img400=8'd33;img401=8'd69;img402=8'd127;img403=8'd116;img404=8'd69;img405=8'd69;img406=8'd69;img407=8'd22;img408=8'd127;img409=8'd127;img410=8'd81;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd17;img436=8'd127;img437=8'd103;img438=8'd11;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd80;img464=8'd127;img465=8'd35;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd43;img491=8'd127;img492=8'd121;img493=8'd25;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd79;img519=8'd127;img520=8'd83;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd116;img547=8'd122;img548=8'd25;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd52;img574=8'd127;img575=8'd116;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd104;img602=8'd127;img603=8'd79;img604=8'd0;img605=8'd7;img606=8'd15;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd104;img630=8'd127;img631=8'd77;img632=8'd46;img633=8'd102;img634=8'd81;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd104;img658=8'd127;img659=8'd127;img660=8'd127;img661=8'd77;img662=8'd15;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd31;img686=8'd95;img687=8'd64;img688=8'd12;img689=8'd3;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd7;img180=8'd75;img181=8'd97;img182=8'd3;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd46;img207=8'd112;img208=8'd127;img209=8'd127;img210=8'd10;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd14;img234=8'd118;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd83;img239=8'd9;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd72;img262=8'd127;img263=8'd127;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd119;img268=8'd58;img269=8'd3;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd16;img289=8'd121;img290=8'd127;img291=8'd104;img292=8'd93;img293=8'd127;img294=8'd127;img295=8'd127;img296=8'd116;img297=8'd12;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd40;img317=8'd127;img318=8'd97;img319=8'd0;img320=8'd4;img321=8'd49;img322=8'd110;img323=8'd127;img324=8'd128;img325=8'd101;img326=8'd9;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd43;img345=8'd127;img346=8'd40;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd91;img351=8'd127;img352=8'd127;img353=8'd96;img354=8'd6;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd88;img373=8'd127;img374=8'd78;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd117;img379=8'd127;img380=8'd127;img381=8'd68;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd43;img401=8'd127;img402=8'd104;img403=8'd20;img404=8'd43;img405=8'd83;img406=8'd126;img407=8'd119;img408=8'd127;img409=8'd118;img410=8'd21;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd9;img429=8'd119;img430=8'd127;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd93;img435=8'd18;img436=8'd108;img437=8'd127;img438=8'd76;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd34;img458=8'd120;img459=8'd128;img460=8'd127;img461=8'd73;img462=8'd4;img463=8'd0;img464=8'd67;img465=8'd127;img466=8'd112;img467=8'd18;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd34;img487=8'd79;img488=8'd71;img489=8'd6;img490=8'd0;img491=8'd0;img492=8'd5;img493=8'd88;img494=8'd127;img495=8'd81;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd44;img522=8'd127;img523=8'd113;img524=8'd9;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd1;img550=8'd83;img551=8'd127;img552=8'd63;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd24;img579=8'd123;img580=8'd127;img581=8'd19;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd58;img608=8'd127;img609=8'd86;img610=8'd5;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd11;img636=8'd109;img637=8'd127;img638=8'd23;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd15;img665=8'd127;img666=8'd83;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd93;img694=8'd122;img695=8'd21;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd7;img722=8'd112;img723=8'd39;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd9;img130=8'd24;img131=8'd24;img132=8'd24;img133=8'd8;img134=8'd65;img135=8'd43;img136=8'd24;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd38;img156=8'd77;img157=8'd109;img158=8'd127;img159=8'd127;img160=8'd127;img161=8'd108;img162=8'd123;img163=8'd127;img164=8'd127;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd18;img181=8'd71;img182=8'd122;img183=8'd126;img184=8'd127;img185=8'd127;img186=8'd127;img187=8'd127;img188=8'd127;img189=8'd127;img190=8'd127;img191=8'd127;img192=8'd127;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd32;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd127;img216=8'd107;img217=8'd85;img218=8'd85;img219=8'd85;img220=8'd85;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd10;img233=8'd66;img234=8'd36;img235=8'd0;img236=8'd29;img237=8'd119;img238=8'd114;img239=8'd119;img240=8'd84;img241=8'd62;img242=8'd35;img243=8'd10;img244=8'd6;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd6;img260=8'd103;img261=8'd127;img262=8'd39;img263=8'd0;img264=8'd0;img265=8'd16;img266=8'd0;img267=8'd15;img268=8'd1;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd3;img287=8'd89;img288=8'd127;img289=8'd66;img290=8'd5;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd6;img314=8'd67;img315=8'd127;img316=8'd117;img317=8'd8;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd46;img342=8'd127;img343=8'd112;img344=8'd14;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd75;img370=8'd127;img371=8'd87;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd117;img398=8'd127;img399=8'd123;img400=8'd64;img401=8'd25;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd128;img426=8'd127;img427=8'd127;img428=8'd127;img429=8'd126;img430=8'd74;img431=8'd46;img432=8'd61;img433=8'd43;img434=8'd21;img435=8'd21;img436=8'd43;img437=8'd14;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd70;img454=8'd127;img455=8'd127;img456=8'd127;img457=8'd127;img458=8'd127;img459=8'd127;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd116;img466=8'd84;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd2;img482=8'd27;img483=8'd109;img484=8'd111;img485=8'd126;img486=8'd127;img487=8'd127;img488=8'd127;img489=8'd127;img490=8'd127;img491=8'd127;img492=8'd127;img493=8'd127;img494=8'd126;img495=8'd62;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd34;img514=8'd36;img515=8'd100;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd127;img520=8'd127;img521=8'd127;img522=8'd127;img523=8'd88;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd60;img544=8'd127;img545=8'd125;img546=8'd76;img547=8'd26;img548=8'd82;img549=8'd127;img550=8'd127;img551=8'd88;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd25;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd94;img576=8'd126;img577=8'd127;img578=8'd127;img579=8'd74;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd5;img600=8'd84;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd125;img606=8'd88;img607=8'd6;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd12;img629=8'd90;img630=8'd116;img631=8'd127;img632=8'd111;img633=8'd64;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd47;img659=8'd75;img660=8'd11;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd18;img210=8'd28;img211=8'd69;img212=8'd101;img213=8'd100;img214=8'd48;img215=8'd19;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd23;img236=8'd76;img237=8'd117;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd127;img243=8'd125;img244=8'd106;img245=8'd76;img246=8'd3;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd23;img262=8'd77;img263=8'd120;img264=8'd127;img265=8'd127;img266=8'd114;img267=8'd83;img268=8'd67;img269=8'd126;img270=8'd100;img271=8'd127;img272=8'd115;img273=8'd113;img274=8'd52;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd77;img289=8'd117;img290=8'd127;img291=8'd127;img292=8'd94;img293=8'd71;img294=8'd4;img295=8'd0;img296=8'd0;img297=8'd96;img298=8'd20;img299=8'd99;img300=8'd123;img301=8'd112;img302=8'd127;img303=8'd11;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd4;img315=8'd63;img316=8'd127;img317=8'd127;img318=8'd117;img319=8'd64;img320=8'd6;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd105;img326=8'd22;img327=8'd35;img328=8'd127;img329=8'd127;img330=8'd127;img331=8'd11;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd36;img343=8'd122;img344=8'd127;img345=8'd114;img346=8'd27;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd2;img352=8'd16;img353=8'd58;img354=8'd113;img355=8'd121;img356=8'd127;img357=8'd128;img358=8'd81;img359=8'd3;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd38;img371=8'd120;img372=8'd127;img373=8'd112;img374=8'd55;img375=8'd69;img376=8'd89;img377=8'd89;img378=8'd85;img379=8'd105;img380=8'd126;img381=8'd116;img382=8'd127;img383=8'd127;img384=8'd127;img385=8'd116;img386=8'd19;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd5;img399=8'd88;img400=8'd122;img401=8'd127;img402=8'd128;img403=8'd127;img404=8'd127;img405=8'd126;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd126;img412=8'd86;img413=8'd13;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd8;img429=8'd68;img430=8'd98;img431=8'd88;img432=8'd73;img433=8'd77;img434=8'd100;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd75;img440=8'd8;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd81;img463=8'd127;img464=8'd127;img465=8'd121;img466=8'd50;img467=8'd2;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd59;img490=8'd125;img491=8'd127;img492=8'd127;img493=8'd45;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd50;img517=8'd121;img518=8'd127;img519=8'd127;img520=8'd106;img521=8'd4;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd27;img544=8'd121;img545=8'd127;img546=8'd127;img547=8'd121;img548=8'd30;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd66;img572=8'd127;img573=8'd127;img574=8'd122;img575=8'd32;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd7;img599=8'd125;img600=8'd127;img601=8'd127;img602=8'd76;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd6;img626=8'd114;img627=8'd127;img628=8'd127;img629=8'd104;img630=8'd4;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd39;img654=8'd128;img655=8'd127;img656=8'd127;img657=8'd33;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd105;img682=8'd127;img683=8'd127;img684=8'd69;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd114;img710=8'd128;img711=8'd117;img712=8'd13;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd57;img738=8'd128;img739=8'd54;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd31;img124=8'd2;img125=8'd21;img126=8'd59;img127=8'd97;img128=8'd59;img129=8'd59;img130=8'd31;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd7;img150=8'd90;img151=8'd123;img152=8'd118;img153=8'd121;img154=8'd127;img155=8'd127;img156=8'd127;img157=8'd127;img158=8'd123;img159=8'd118;img160=8'd42;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd76;img178=8'd127;img179=8'd127;img180=8'd127;img181=8'd107;img182=8'd96;img183=8'd89;img184=8'd89;img185=8'd90;img186=8'd127;img187=8'd127;img188=8'd121;img189=8'd23;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd22;img205=8'd118;img206=8'd127;img207=8'd113;img208=8'd32;img209=8'd14;img210=8'd6;img211=8'd0;img212=8'd0;img213=8'd1;img214=8'd64;img215=8'd126;img216=8'd128;img217=8'd87;img218=8'd9;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd28;img233=8'd127;img234=8'd127;img235=8'd54;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd67;img244=8'd125;img245=8'd127;img246=8'd38;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd32;img261=8'd127;img262=8'd79;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd111;img273=8'd127;img274=8'd79;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd97;img289=8'd127;img290=8'd52;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd75;img301=8'd127;img302=8'd107;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd17;img316=8'd110;img317=8'd120;img318=8'd29;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd42;img329=8'd127;img330=8'd107;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd63;img344=8'd127;img345=8'd86;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd42;img357=8'd127;img358=8'd107;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd107;img372=8'd120;img373=8'd30;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd42;img385=8'd127;img386=8'd107;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd107;img400=8'd100;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd42;img413=8'd127;img414=8'd107;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd6;img427=8'd110;img428=8'd100;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd42;img441=8'd127;img442=8'd107;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd49;img455=8'd127;img456=8'd100;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd81;img469=8'd127;img470=8'd105;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd49;img483=8'd127;img484=8'd100;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd26;img496=8'd119;img497=8'd127;img498=8'd38;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd49;img511=8'd127;img512=8'd100;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd26;img523=8'd83;img524=8'd127;img525=8'd98;img526=8'd2;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd33;img539=8'd121;img540=8'd100;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd2;img550=8'd84;img551=8'd127;img552=8'd114;img553=8'd28;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd107;img568=8'd107;img569=8'd10;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd23;img576=8'd76;img577=8'd101;img578=8'd127;img579=8'd127;img580=8'd32;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd107;img596=8'd127;img597=8'd102;img598=8'd90;img599=8'd90;img600=8'd90;img601=8'd90;img602=8'd90;img603=8'd118;img604=8'd127;img605=8'd127;img606=8'd117;img607=8'd78;img608=8'd5;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd41;img624=8'd103;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd127;img629=8'd127;img630=8'd127;img631=8'd127;img632=8'd126;img633=8'd117;img634=8'd60;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd13;img653=8'd105;img654=8'd127;img655=8'd127;img656=8'd127;img657=8'd127;img658=8'd127;img659=8'd77;img660=8'd52;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd4;img95=8'd102;img96=8'd127;img97=8'd88;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd4;img122=8'd75;img123=8'd126;img124=8'd126;img125=8'd63;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd59;img150=8'd126;img151=8'd93;img152=8'd28;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd71;img178=8'd126;img179=8'd59;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd77;img206=8'd124;img207=8'd25;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd13;img233=8'd127;img234=8'd98;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd75;img261=8'd127;img262=8'd98;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd29;img271=8'd43;img272=8'd43;img273=8'd19;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd113;img289=8'd127;img290=8'd48;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd76;img297=8'd113;img298=8'd122;img299=8'd126;img300=8'd126;img301=8'd119;img302=8'd63;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd5;img316=8'd115;img317=8'd113;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd2;img322=8'd27;img323=8'd115;img324=8'd127;img325=8'd128;img326=8'd117;img327=8'd88;img328=8'd113;img329=8'd128;img330=8'd114;img331=8'd16;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd55;img344=8'd126;img345=8'd75;img346=8'd0;img347=8'd0;img348=8'd13;img349=8'd64;img350=8'd126;img351=8'd126;img352=8'd114;img353=8'd67;img354=8'd14;img355=8'd0;img356=8'd0;img357=8'd89;img358=8'd126;img359=8'd28;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd80;img372=8'd126;img373=8'd57;img374=8'd0;img375=8'd0;img376=8'd75;img377=8'd127;img378=8'd126;img379=8'd93;img380=8'd22;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd71;img386=8'd126;img387=8'd28;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd93;img400=8'd126;img401=8'd57;img402=8'd0;img403=8'd19;img404=8'd119;img405=8'd127;img406=8'd76;img407=8'd3;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd71;img414=8'd101;img415=8'd3;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd99;img428=8'd127;img429=8'd57;img430=8'd0;img431=8'd74;img432=8'd127;img433=8'd82;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd77;img442=8'd99;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd99;img456=8'd126;img457=8'd57;img458=8'd0;img459=8'd86;img460=8'd126;img461=8'd94;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd13;img469=8'd127;img470=8'd86;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd99;img484=8'd126;img485=8'd57;img486=8'd0;img487=8'd10;img488=8'd116;img489=8'd124;img490=8'd61;img491=8'd10;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd100;img497=8'd122;img498=8'd28;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd13;img511=8'd111;img512=8'd126;img513=8'd57;img514=8'd0;img515=8'd0;img516=8'd13;img517=8'd102;img518=8'd126;img519=8'd97;img520=8'd7;img521=8'd0;img522=8'd38;img523=8'd100;img524=8'd125;img525=8'd63;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd93;img540=8'd127;img541=8'd90;img542=8'd5;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd38;img547=8'd18;img548=8'd15;img549=8'd77;img550=8'd127;img551=8'd122;img552=8'd63;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd14;img568=8'd105;img569=8'd127;img570=8'd98;img571=8'd41;img572=8'd29;img573=8'd29;img574=8'd66;img575=8'd99;img576=8'd126;img577=8'd127;img578=8'd107;img579=8'd41;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd13;img597=8'd108;img598=8'd126;img599=8'd126;img600=8'd126;img601=8'd127;img602=8'd126;img603=8'd126;img604=8'd126;img605=8'd78;img606=8'd10;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd8;img626=8'd52;img627=8'd70;img628=8'd120;img629=8'd70;img630=8'd70;img631=8'd70;img632=8'd20;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd25;img209=8'd90;img210=8'd127;img211=8'd128;img212=8'd127;img213=8'd85;img214=8'd18;img215=8'd6;img216=8'd38;img217=8'd5;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd3;img235=8'd34;img236=8'd114;img237=8'd126;img238=8'd126;img239=8'd127;img240=8'd126;img241=8'd126;img242=8'd80;img243=8'd95;img244=8'd127;img245=8'd46;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd28;img263=8'd126;img264=8'd126;img265=8'd114;img266=8'd40;img267=8'd35;img268=8'd35;img269=8'd50;img270=8'd45;img271=8'd118;img272=8'd124;img273=8'd34;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd22;img290=8'd117;img291=8'd126;img292=8'd93;img293=8'd25;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd13;img298=8'd102;img299=8'd126;img300=8'd68;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd84;img318=8'd127;img319=8'd89;img320=8'd19;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd35;img326=8'd126;img327=8'd126;img328=8'd32;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd78;img345=8'd127;img346=8'd121;img347=8'd21;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd3;img353=8'd96;img354=8'd127;img355=8'd95;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd104;img373=8'd126;img374=8'd115;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd3;img380=8'd68;img381=8'd126;img382=8'd126;img383=8'd32;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd104;img401=8'd126;img402=8'd115;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd16;img407=8'd69;img408=8'd126;img409=8'd126;img410=8'd114;img411=8'd8;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd83;img429=8'd126;img430=8'd125;img431=8'd104;img432=8'd104;img433=8'd104;img434=8'd114;img435=8'd127;img436=8'd126;img437=8'd126;img438=8'd80;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd5;img457=8'd90;img458=8'd127;img459=8'd126;img460=8'd126;img461=8'd126;img462=8'd126;img463=8'd38;img464=8'd85;img465=8'd126;img466=8'd28;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd32;img487=8'd58;img488=8'd58;img489=8'd37;img490=8'd0;img491=8'd75;img492=8'd127;img493=8'd108;img494=8'd11;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd127;img520=8'd126;img521=8'd81;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd16;img547=8'd127;img548=8'd120;img549=8'd25;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd79;img575=8'd127;img576=8'd82;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd22;img602=8'd120;img603=8'd127;img604=8'd46;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd47;img630=8'd127;img631=8'd126;img632=8'd42;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd57;img658=8'd126;img659=8'd105;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd104;img686=8'd126;img687=8'd58;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd83;img714=8'd126;img715=8'd58;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd47;img742=8'd100;img743=8'd32;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd9;img153=8'd33;img154=8'd69;img155=8'd128;img156=8'd127;img157=8'd85;img158=8'd69;img159=8'd12;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd3;img179=8'd60;img180=8'd114;img181=8'd126;img182=8'd126;img183=8'd127;img184=8'd126;img185=8'd126;img186=8'd126;img187=8'd79;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd54;img207=8'd126;img208=8'd126;img209=8'd126;img210=8'd126;img211=8'd95;img212=8'd126;img213=8'd126;img214=8'd126;img215=8'd126;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd22;img234=8'd117;img235=8'd126;img236=8'd126;img237=8'd126;img238=8'd58;img239=8'd3;img240=8'd68;img241=8'd126;img242=8'd126;img243=8'd126;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd22;img261=8'd89;img262=8'd127;img263=8'd126;img264=8'd111;img265=8'd22;img266=8'd1;img267=8'd0;img268=8'd3;img269=8'd27;img270=8'd116;img271=8'd126;img272=8'd105;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd47;img289=8'd127;img290=8'd128;img291=8'd125;img292=8'd58;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd68;img299=8'd126;img300=8'd128;img301=8'd77;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd83;img317=8'd126;img318=8'd127;img319=8'd93;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd105;img328=8'd127;img329=8'd103;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd10;img344=8'd110;img345=8'd126;img346=8'd127;img347=8'd46;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd58;img356=8'd127;img357=8'd103;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd35;img372=8'd126;img373=8'd126;img374=8'd96;img375=8'd9;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd58;img384=8'd127;img385=8'd112;img386=8'd13;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd61;img400=8'd126;img401=8'd126;img402=8'd32;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd58;img412=8'd127;img413=8'd126;img414=8'd35;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd66;img428=8'd127;img429=8'd127;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd58;img440=8'd128;img441=8'd127;img442=8'd35;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd92;img456=8'd126;img457=8'd126;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd58;img468=8'd127;img469=8'd126;img470=8'd35;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd92;img484=8'd126;img485=8'd126;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd58;img496=8'd127;img497=8'd120;img498=8'd25;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd92;img512=8'd126;img513=8'd126;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd105;img524=8'd127;img525=8'd56;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd24;img540=8'd116;img541=8'd126;img542=8'd79;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd115;img552=8'd116;img553=8'd4;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd47;img569=8'd127;img570=8'd122;img571=8'd25;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd78;img579=8'd127;img580=8'd84;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd17;img597=8'd82;img598=8'd127;img599=8'd57;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd33;img606=8'd118;img607=8'd116;img608=8'd21;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd16;img626=8'd111;img627=8'd120;img628=8'd67;img629=8'd0;img630=8'd0;img631=8'd19;img632=8'd46;img633=8'd117;img634=8'd126;img635=8'd69;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd13;img655=8'd89;img656=8'd120;img657=8'd104;img658=8'd52;img659=8'd117;img660=8'd126;img661=8'd126;img662=8'd88;img663=8'd18;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd8;img684=8'd27;img685=8'd90;img686=8'd126;img687=8'd69;img688=8'd69;img689=8'd27;img690=8'd2;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd64;img126=8'd128;img127=8'd96;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd96;img154=8'd128;img155=8'd128;img156=8'd32;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd128;img182=8'd128;img183=8'd128;img184=8'd64;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd128;img210=8'd128;img211=8'd128;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd128;img238=8'd128;img239=8'd128;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd64;img266=8'd128;img267=8'd128;img268=8'd64;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd128;img294=8'd128;img295=8'd128;img296=8'd64;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd128;img322=8'd128;img323=8'd128;img324=8'd64;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd128;img350=8'd128;img351=8'd128;img352=8'd64;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd128;img378=8'd128;img379=8'd128;img380=8'd64;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd128;img406=8'd128;img407=8'd128;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd128;img434=8'd128;img435=8'd128;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd128;img462=8'd128;img463=8'd128;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd128;img490=8'd128;img491=8'd128;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd96;img518=8'd128;img519=8'd128;img520=8'd64;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd96;img546=8'd128;img547=8'd128;img548=8'd64;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd32;img573=8'd128;img574=8'd128;img575=8'd128;img576=8'd64;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd96;img601=8'd128;img602=8'd128;img603=8'd128;img604=8'd64;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd32;img628=8'd128;img629=8'd128;img630=8'd128;img631=8'd32;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd32;img656=8'd128;img657=8'd64;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd26;img125=8'd66;img126=8'd107;img127=8'd127;img128=8'd127;img129=8'd127;img130=8'd102;img131=8'd81;img132=8'd21;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd51;img149=8'd71;img150=8'd102;img151=8'd102;img152=8'd127;img153=8'd126;img154=8'd127;img155=8'd126;img156=8'd76;img157=8'd35;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd127;img177=8'd127;img178=8'd122;img179=8'd102;img180=8'd71;img181=8'd51;img182=8'd41;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd86;img205=8'd126;img206=8'd102;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd11;img233=8'd112;img234=8'd117;img235=8'd15;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd61;img262=8'd127;img263=8'd25;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd62;img290=8'd127;img291=8'd46;img292=8'd26;img293=8'd26;img294=8'd26;img295=8'd5;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd11;img317=8'd112;img318=8'd127;img319=8'd126;img320=8'd127;img321=8'd126;img322=8'd127;img323=8'd86;img324=8'd41;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd11;img344=8'd107;img345=8'd127;img346=8'd102;img347=8'd81;img348=8'd51;img349=8'd51;img350=8'd102;img351=8'd112;img352=8'd127;img353=8'd127;img354=8'd26;img355=8'd5;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd31;img372=8'd127;img373=8'd86;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd10;img380=8'd56;img381=8'd96;img382=8'd127;img383=8'd106;img384=8'd21;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd51;img411=8'd102;img412=8'd117;img413=8'd26;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd10;img440=8'd107;img441=8'd116;img442=8'd41;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd31;img469=8'd102;img470=8'd117;img471=8'd56;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd10;img498=8'd107;img499=8'd126;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd77;img527=8'd127;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd21;img554=8'd117;img555=8'd106;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd57;img569=8'd46;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd16;img581=8'd87;img582=8'd122;img583=8'd20;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd41;img596=8'd127;img597=8'd76;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd11;img605=8'd51;img606=8'd51;img607=8'd92;img608=8'd117;img609=8'd106;img610=8'd41;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd41;img624=8'd128;img625=8'd127;img626=8'd117;img627=8'd76;img628=8'd77;img629=8'd97;img630=8'd87;img631=8'd127;img632=8'd127;img633=8'd127;img634=8'd127;img635=8'd107;img636=8'd71;img637=8'd10;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd36;img653=8'd76;img654=8'd76;img655=8'd116;img656=8'd127;img657=8'd106;img658=8'd96;img659=8'd76;img660=8'd66;img661=8'd25;img662=8'd25;img663=8'd5;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd32;img180=8'd73;img181=8'd115;img182=8'd128;img183=8'd103;img184=8'd60;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd12;img206=8'd99;img207=8'd126;img208=8'd127;img209=8'd113;img210=8'd108;img211=8'd118;img212=8'd126;img213=8'd45;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd10;img233=8'd103;img234=8'd127;img235=8'd112;img236=8'd35;img237=8'd8;img238=8'd0;img239=8'd15;img240=8'd103;img241=8'd87;img242=8'd1;img243=8'd44;img244=8'd19;img245=8'd1;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd69;img261=8'd127;img262=8'd114;img263=8'd3;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd18;img269=8'd14;img270=8'd38;img271=8'd127;img272=8'd127;img273=8'd5;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd44;img288=8'd126;img289=8'd118;img290=8'd6;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd21;img298=8'd119;img299=8'd127;img300=8'd87;img301=8'd1;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd67;img316=8'd127;img317=8'd96;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd7;img326=8'd119;img327=8'd127;img328=8'd81;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd85;img344=8'd127;img345=8'd37;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd43;img354=8'd124;img355=8'd127;img356=8'd38;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd5;img371=8'd125;img372=8'd127;img373=8'd24;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd3;img381=8'd110;img382=8'd127;img383=8'd121;img384=8'd16;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd5;img399=8'd127;img400=8'd127;img401=8'd24;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd3;img408=8'd36;img409=8'd127;img410=8'd127;img411=8'd72;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd3;img427=8'd111;img428=8'd127;img429=8'd59;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd13;img435=8'd59;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd24;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd14;img456=8'd121;img457=8'd127;img458=8'd94;img459=8'd52;img460=8'd73;img461=8'd80;img462=8'd110;img463=8'd122;img464=8'd120;img465=8'd127;img466=8'd112;img467=8'd9;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd39;img485=8'd101;img486=8'd127;img487=8'd127;img488=8'd124;img489=8'd108;img490=8'd78;img491=8'd34;img492=8'd124;img493=8'd127;img494=8'd79;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd3;img514=8'd28;img515=8'd28;img516=8'd25;img517=8'd0;img518=8'd0;img519=8'd19;img520=8'd127;img521=8'd127;img522=8'd37;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd33;img548=8'd127;img549=8'd127;img550=8'd9;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd75;img576=8'd127;img577=8'd127;img578=8'd9;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd15;img603=8'd119;img604=8'd127;img605=8'd96;img606=8'd2;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd33;img631=8'd127;img632=8'd127;img633=8'd56;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd44;img659=8'd127;img660=8'd122;img661=8'd2;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd85;img687=8'd127;img688=8'd99;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd127;img715=8'd127;img716=8'd75;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd37;img201=8'd125;img202=8'd127;img203=8'd127;img204=8'd127;img205=8'd123;img206=8'd84;img207=8'd84;img208=8'd68;img209=8'd13;img210=8'd40;img211=8'd30;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd52;img229=8'd127;img230=8'd127;img231=8'd127;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd125;img238=8'd127;img239=8'd126;img240=8'd99;img241=8'd57;img242=8'd36;img243=8'd20;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd3;img257=8'd50;img258=8'd68;img259=8'd53;img260=8'd53;img261=8'd57;img262=8'd96;img263=8'd96;img264=8'd96;img265=8'd117;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd127;img270=8'd127;img271=8'd123;img272=8'd65;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd23;img294=8'd57;img295=8'd57;img296=8'd102;img297=8'd127;img298=8'd127;img299=8'd127;img300=8'd120;img301=8'd8;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd4;img325=8'd18;img326=8'd78;img327=8'd127;img328=8'd127;img329=8'd65;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd18;img355=8'd127;img356=8'd121;img357=8'd17;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd58;img383=8'd127;img384=8'd127;img385=8'd59;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd17;img410=8'd122;img411=8'd127;img412=8'd120;img413=8'd9;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd56;img438=8'd127;img439=8'd127;img440=8'd70;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd19;img465=8'd122;img466=8'd127;img467=8'd122;img468=8'd20;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd10;img492=8'd88;img493=8'd127;img494=8'd127;img495=8'd57;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd70;img520=8'd127;img521=8'd127;img522=8'd110;img523=8'd1;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd44;img547=8'd127;img548=8'd127;img549=8'd122;img550=8'd23;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd32;img574=8'd121;img575=8'd127;img576=8'd127;img577=8'd42;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd8;img601=8'd122;img602=8'd127;img603=8'd127;img604=8'd74;img605=8'd3;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd1;img628=8'd56;img629=8'd127;img630=8'd127;img631=8'd102;img632=8'd3;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd29;img656=8'd127;img657=8'd127;img658=8'd127;img659=8'd42;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd7;img683=8'd119;img684=8'd127;img685=8'd128;img686=8'd97;img687=8'd2;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd41;img711=8'd127;img712=8'd127;img713=8'd97;img714=8'd14;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd20;img739=8'd115;img740=8'd97;img741=8'd14;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd6;img119=8'd21;img120=8'd73;img121=8'd73;img122=8'd24;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd6;img146=8'd65;img147=8'd127;img148=8'd127;img149=8'd127;img150=8'd125;img151=8'd82;img152=8'd9;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd67;img174=8'd127;img175=8'd127;img176=8'd127;img177=8'd127;img178=8'd127;img179=8'd127;img180=8'd115;img181=8'd35;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd51;img202=8'd127;img203=8'd126;img204=8'd73;img205=8'd51;img206=8'd54;img207=8'd119;img208=8'd127;img209=8'd124;img210=8'd64;img211=8'd5;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd91;img230=8'd127;img231=8'd84;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd31;img236=8'd118;img237=8'd127;img238=8'd127;img239=8'd82;img240=8'd3;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd128;img258=8'd127;img259=8'd22;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd29;img265=8'd97;img266=8'd127;img267=8'd127;img268=8'd82;img269=8'd2;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd94;img286=8'd127;img287=8'd16;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd28;img294=8'd118;img295=8'd127;img296=8'd127;img297=8'd43;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd73;img314=8'd127;img315=8'd16;img316=8'd0;img317=8'd50;img318=8'd95;img319=8'd44;img320=8'd44;img321=8'd44;img322=8'd74;img323=8'd127;img324=8'd127;img325=8'd62;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd47;img342=8'd127;img343=8'd39;img344=8'd20;img345=8'd124;img346=8'd127;img347=8'd127;img348=8'd127;img349=8'd127;img350=8'd127;img351=8'd127;img352=8'd127;img353=8'd112;img354=8'd42;img355=8'd8;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd7;img370=8'd46;img371=8'd6;img372=8'd18;img373=8'd120;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd127;img383=8'd122;img384=8'd45;img385=8'd5;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd38;img402=8'd81;img403=8'd90;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd127;img413=8'd105;img414=8'd22;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd2;img432=8'd8;img433=8'd8;img434=8'd20;img435=8'd19;img436=8'd8;img437=8'd8;img438=8'd73;img439=8'd122;img440=8'd127;img441=8'd127;img442=8'd93;img443=8'd24;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd10;img458=8'd29;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd29;img468=8'd105;img469=8'd127;img470=8'd127;img471=8'd92;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd39;img485=8'd111;img486=8'd124;img487=8'd40;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd7;img497=8'd110;img498=8'd127;img499=8'd120;img500=8'd36;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd45;img513=8'd124;img514=8'd127;img515=8'd126;img516=8'd29;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd27;img526=8'd126;img527=8'd127;img528=8'd96;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd58;img542=8'd127;img543=8'd127;img544=8'd30;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd50;img554=8'd126;img555=8'd127;img556=8'd73;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd7;img570=8'd94;img571=8'd127;img572=8'd111;img573=8'd79;img574=8'd19;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd56;img580=8'd106;img581=8'd123;img582=8'd127;img583=8'd127;img584=8'd73;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd6;img599=8'd111;img600=8'd123;img601=8'd127;img602=8'd126;img603=8'd125;img604=8'd125;img605=8'd125;img606=8'd125;img607=8'd127;img608=8'd127;img609=8'd127;img610=8'd127;img611=8'd100;img612=8'd10;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd48;img629=8'd92;img630=8'd114;img631=8'd127;img632=8'd127;img633=8'd127;img634=8'd127;img635=8'd127;img636=8'd127;img637=8'd98;img638=8'd62;img639=8'd12;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd12;img659=8'd19;img660=8'd69;img661=8'd37;img662=8'd63;img663=8'd44;img664=8'd19;img665=8'd4;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd84;img159=8'd46;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd1;img186=8'd117;img187=8'd63;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd26;img214=8'd127;img215=8'd63;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd19;img234=8'd89;img235=8'd16;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd26;img242=8'd127;img243=8'd41;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd47;img262=8'd127;img263=8'd42;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd44;img270=8'd127;img271=8'd27;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd80;img290=8'd127;img291=8'd28;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd95;img298=8'd119;img299=8'd2;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd7;img317=8'd114;img318=8'd84;img319=8'd1;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd97;img326=8'd118;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd28;img345=8'd127;img346=8'd57;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd8;img353=8'd118;img354=8'd84;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd58;img373=8'd127;img374=8'd25;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd52;img381=8'd127;img382=8'd53;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd4;img400=8'd111;img401=8'd118;img402=8'd38;img403=8'd78;img404=8'd90;img405=8'd95;img406=8'd126;img407=8'd126;img408=8'd127;img409=8'd127;img410=8'd57;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd8;img428=8'd127;img429=8'd127;img430=8'd127;img431=8'd126;img432=8'd106;img433=8'd90;img434=8'd90;img435=8'd90;img436=8'd123;img437=8'd127;img438=8'd124;img439=8'd47;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd4;img456=8'd109;img457=8'd120;img458=8'd59;img459=8'd11;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd113;img465=8'd127;img466=8'd121;img467=8'd99;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd7;img485=8'd9;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd14;img492=8'd122;img493=8'd104;img494=8'd23;img495=8'd19;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd50;img520=8'd127;img521=8'd66;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd58;img548=8'd127;img549=8'd34;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd58;img576=8'd127;img577=8'd31;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd58;img604=8'd127;img605=8'd31;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd87;img632=8'd128;img633=8'd50;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd94;img660=8'd127;img661=8'd42;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd58;img688=8'd88;img689=8'd5;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd16;img184=8'd70;img185=8'd97;img186=8'd22;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd19;img210=8'd73;img211=8'd120;img212=8'd127;img213=8'd127;img214=8'd114;img215=8'd24;img216=8'd39;img217=8'd23;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd1;img236=8'd22;img237=8'd115;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd127;img243=8'd121;img244=8'd127;img245=8'd99;img246=8'd1;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd11;img263=8'd65;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd120;img268=8'd126;img269=8'd127;img270=8'd127;img271=8'd127;img272=8'd127;img273=8'd119;img274=8'd2;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd77;img291=8'd127;img292=8'd127;img293=8'd125;img294=8'd52;img295=8'd36;img296=8'd99;img297=8'd127;img298=8'd127;img299=8'd127;img300=8'd117;img301=8'd29;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd1;img317=8'd87;img318=8'd126;img319=8'd126;img320=8'd103;img321=8'd26;img322=8'd60;img323=8'd108;img324=8'd127;img325=8'd127;img326=8'd127;img327=8'd127;img328=8'd92;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd56;img345=8'd127;img346=8'd127;img347=8'd108;img348=8'd44;img349=8'd124;img350=8'd127;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd127;img355=8'd109;img356=8'd16;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd3;img372=8'd116;img373=8'd127;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd118;img379=8'd64;img380=8'd98;img381=8'd127;img382=8'd127;img383=8'd60;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd2;img400=8'd99;img401=8'd127;img402=8'd127;img403=8'd123;img404=8'd119;img405=8'd66;img406=8'd9;img407=8'd23;img408=8'd124;img409=8'd127;img410=8'd100;img411=8'd7;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd8;img429=8'd46;img430=8'd44;img431=8'd20;img432=8'd0;img433=8'd0;img434=8'd6;img435=8'd87;img436=8'd127;img437=8'd121;img438=8'd19;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd48;img463=8'd127;img464=8'd127;img465=8'd78;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd9;img490=8'd105;img491=8'd127;img492=8'd113;img493=8'd3;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd99;img518=8'd127;img519=8'd127;img520=8'd50;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd17;img545=8'd121;img546=8'd127;img547=8'd90;img548=8'd2;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd14;img572=8'd112;img573=8'd127;img574=8'd113;img575=8'd15;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd39;img600=8'd127;img601=8'd128;img602=8'd64;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd27;img627=8'd119;img628=8'd127;img629=8'd124;img630=8'd27;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd6;img654=8'd92;img655=8'd127;img656=8'd127;img657=8'd116;img658=8'd21;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd57;img682=8'd127;img683=8'd127;img684=8'd115;img685=8'd24;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd55;img710=8'd120;img711=8'd63;img712=8'd13;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd25;img97=8'd90;img98=8'd127;img99=8'd122;img100=8'd25;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd92;img125=8'd126;img126=8'd126;img127=8'd116;img128=8'd82;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd33;img152=8'd117;img153=8'd126;img154=8'd68;img155=8'd19;img156=8'd28;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd10;img179=8'd118;img180=8'd126;img181=8'd88;img182=8'd2;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd38;img207=8'd126;img208=8'd126;img209=8'd28;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd70;img235=8'd127;img236=8'd87;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd11;img262=8'd106;img263=8'd126;img264=8'd35;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd58;img290=8'd127;img291=8'd120;img292=8'd25;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd79;img318=8'd127;img319=8'd103;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd115;img346=8'd127;img347=8'd51;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd116;img374=8'd128;img375=8'd90;img376=8'd69;img377=8'd90;img378=8'd127;img379=8'd128;img380=8'd127;img381=8'd111;img382=8'd49;img383=8'd2;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd115;img402=8'd127;img403=8'd126;img404=8'd126;img405=8'd126;img406=8'd126;img407=8'd106;img408=8'd126;img409=8'd126;img410=8'd126;img411=8'd59;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd115;img430=8'd127;img431=8'd120;img432=8'd92;img433=8'd45;img434=8'd35;img435=8'd4;img436=8'd35;img437=8'd86;img438=8'd126;img439=8'd126;img440=8'd43;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd68;img458=8'd127;img459=8'd77;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd7;img466=8'd108;img467=8'd126;img468=8'd58;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd58;img486=8'd127;img487=8'd103;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd78;img495=8'd126;img496=8'd58;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd53;img514=8'd128;img515=8'd106;img516=8'd4;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd25;img522=8'd117;img523=8'd127;img524=8'd58;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd80;img543=8'd126;img544=8'd77;img545=8'd5;img546=8'd0;img547=8'd0;img548=8'd15;img549=8'd99;img550=8'd126;img551=8'd126;img552=8'd48;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd9;img571=8'd114;img572=8'd126;img573=8'd77;img574=8'd35;img575=8'd41;img576=8'd114;img577=8'd126;img578=8'd114;img579=8'd65;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd25;img600=8'd114;img601=8'd126;img602=8'd126;img603=8'd127;img604=8'd126;img605=8'd93;img606=8'd25;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd24;img629=8'd90;img630=8'd126;img631=8'd95;img632=8'd59;img633=8'd3;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd57;img94=8'd128;img95=8'd29;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd113;img122=8'd128;img123=8'd29;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd15;img149=8'd128;img150=8'd57;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd57;img177=8'd128;img178=8'd43;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd99;img205=8'd128;img206=8'd15;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd15;img232=8'd128;img233=8'd113;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd71;img260=8'd128;img261=8'd71;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd29;img269=8'd43;img270=8'd43;img271=8'd71;img272=8'd29;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd85;img288=8'd128;img289=8'd43;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd29;img296=8'd113;img297=8'd128;img298=8'd128;img299=8'd128;img300=8'd128;img301=8'd29;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd85;img316=8'd128;img317=8'd43;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd85;img324=8'd128;img325=8'd128;img326=8'd57;img327=8'd29;img328=8'd113;img329=8'd99;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd85;img344=8'd128;img345=8'd43;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd29;img351=8'd128;img352=8'd128;img353=8'd43;img354=8'd0;img355=8'd0;img356=8'd85;img357=8'd128;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd85;img372=8'd128;img373=8'd43;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd85;img379=8'd128;img380=8'd43;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd85;img385=8'd128;img386=8'd43;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd71;img400=8'd128;img401=8'd57;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd15;img406=8'd128;img407=8'd99;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd85;img413=8'd128;img414=8'd43;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd15;img428=8'd128;img429=8'd128;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd85;img434=8'd128;img435=8'd57;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd99;img441=8'd113;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd99;img457=8'd128;img458=8'd57;img459=8'd0;img460=8'd0;img461=8'd85;img462=8'd128;img463=8'd43;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd43;img468=8'd128;img469=8'd57;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd43;img485=8'd128;img486=8'd128;img487=8'd85;img488=8'd29;img489=8'd128;img490=8'd128;img491=8'd15;img492=8'd0;img493=8'd0;img494=8'd43;img495=8'd113;img496=8'd113;img497=8'd15;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd57;img514=8'd113;img515=8'd128;img516=8'd128;img517=8'd128;img518=8'd128;img519=8'd43;img520=8'd43;img521=8'd85;img522=8'd128;img523=8'd128;img524=8'd29;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd15;img543=8'd71;img544=8'd128;img545=8'd128;img546=8'd128;img547=8'd128;img548=8'd128;img549=8'd128;img550=8'd99;img551=8'd15;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd113;img574=8'd128;img575=8'd128;img576=8'd71;img577=8'd43;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd71;img602=8'd128;img603=8'd128;img604=8'd85;img605=8'd85;img606=8'd29;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd71;img631=8'd113;img632=8'd85;img633=8'd57;img634=8'd15;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd35;img157=8'd76;img158=8'd119;img159=8'd127;img160=8'd127;img161=8'd128;img162=8'd127;img163=8'd126;img164=8'd26;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd44;img182=8'd82;img183=8'd119;img184=8'd127;img185=8'd127;img186=8'd109;img187=8'd69;img188=8'd42;img189=8'd20;img190=8'd77;img191=8'd127;img192=8'd68;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd69;img208=8'd123;img209=8'd127;img210=8'd127;img211=8'd108;img212=8'd84;img213=8'd27;img214=8'd3;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd50;img219=8'd96;img220=8'd2;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd117;img236=8'd127;img237=8'd85;img238=8'd27;img239=8'd3;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd18;img247=8'd4;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd87;img264=8'd127;img265=8'd47;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd19;img291=8'd123;img292=8'd111;img293=8'd7;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd71;img319=8'd127;img320=8'd75;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd76;img347=8'd127;img348=8'd56;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd113;img375=8'd121;img376=8'd16;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd6;img402=8'd120;img403=8'd102;img404=8'd22;img405=8'd22;img406=8'd22;img407=8'd22;img408=8'd4;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd35;img430=8'd127;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd103;img437=8'd43;img438=8'd4;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd19;img458=8'd92;img459=8'd85;img460=8'd67;img461=8'd67;img462=8'd81;img463=8'd106;img464=8'd127;img465=8'd127;img466=8'd83;img467=8'd4;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd5;img492=8'd26;img493=8'd89;img494=8'd127;img495=8'd63;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd14;img521=8'd105;img522=8'd127;img523=8'd52;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd32;img548=8'd105;img549=8'd127;img550=8'd97;img551=8'd7;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd3;img572=8'd0;img573=8'd5;img574=8'd69;img575=8'd122;img576=8'd127;img577=8'd99;img578=8'd26;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd7;img598=8'd44;img599=8'd61;img600=8'd74;img601=8'd112;img602=8'd127;img603=8'd124;img604=8'd64;img605=8'd7;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd2;img624=8'd59;img625=8'd125;img626=8'd105;img627=8'd124;img628=8'd127;img629=8'd126;img630=8'd100;img631=8'd25;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd69;img652=8'd127;img653=8'd127;img654=8'd127;img655=8'd125;img656=8'd101;img657=8'd36;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd40;img680=8'd84;img681=8'd99;img682=8'd44;img683=8'd4;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd99;img152=8'd30;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd25;img179=8'd122;img180=8'd21;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd1;img206=8'd93;img207=8'd118;img208=8'd11;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd67;img213=8'd42;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd44;img234=8'd107;img235=8'd13;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd65;img241=8'd85;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd64;img262=8'd60;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd46;img269=8'd105;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd16;img289=8'd117;img290=8'd56;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd46;img297=8'd121;img298=8'd15;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd58;img317=8'd111;img318=8'd11;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd85;img325=8'd122;img326=8'd29;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd15;img344=8'd120;img345=8'd62;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd20;img352=8'd125;img353=8'd69;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd2;img371=8'd64;img372=8'd121;img373=8'd9;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd8;img380=8'd115;img381=8'd67;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd8;img399=8'd127;img400=8'd90;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd83;img409=8'd67;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd5;img427=8'd96;img428=8'd117;img429=8'd68;img430=8'd51;img431=8'd10;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd57;img437=8'd108;img438=8'd16;img439=8'd16;img440=8'd16;img441=8'd1;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd4;img456=8'd45;img457=8'd64;img458=8'd97;img459=8'd109;img460=8'd105;img461=8'd105;img462=8'd106;img463=8'd105;img464=8'd113;img465=8'd127;img466=8'd127;img467=8'd102;img468=8'd60;img469=8'd4;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd5;img488=8'd8;img489=8'd19;img490=8'd45;img491=8'd45;img492=8'd98;img493=8'd121;img494=8'd17;img495=8'd3;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd83;img521=8'd117;img522=8'd8;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd83;img549=8'd72;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd46;img577=8'd94;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd46;img605=8'd117;img606=8'd17;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd10;img633=8'd127;img634=8'd31;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd2;img661=8'd105;img662=8'd110;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd54;img690=8'd83;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd2;img126=8'd40;img127=8'd98;img128=8'd43;img129=8'd40;img130=8'd40;img131=8'd40;img132=8'd7;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd5;img154=8'd127;img155=8'd127;img156=8'd127;img157=8'd127;img158=8'd127;img159=8'd127;img160=8'd76;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd6;img178=8'd31;img179=8'd28;img180=8'd0;img181=8'd5;img182=8'd127;img183=8'd127;img184=8'd127;img185=8'd127;img186=8'd127;img187=8'd127;img188=8'd126;img189=8'd119;img190=8'd29;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd71;img206=8'd127;img207=8'd121;img208=8'd42;img209=8'd2;img210=8'd81;img211=8'd127;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd127;img216=8'd127;img217=8'd127;img218=8'd30;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd6;img232=8'd71;img233=8'd124;img234=8'd127;img235=8'd127;img236=8'd74;img237=8'd0;img238=8'd37;img239=8'd105;img240=8'd126;img241=8'd127;img242=8'd127;img243=8'd127;img244=8'd127;img245=8'd127;img246=8'd106;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd74;img260=8'd127;img261=8'd127;img262=8'd127;img263=8'd127;img264=8'd100;img265=8'd17;img266=8'd0;img267=8'd0;img268=8'd80;img269=8'd127;img270=8'd71;img271=8'd97;img272=8'd127;img273=8'd127;img274=8'd122;img275=8'd39;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd5;img286=8'd68;img287=8'd125;img288=8'd127;img289=8'd127;img290=8'd127;img291=8'd127;img292=8'd127;img293=8'd35;img294=8'd0;img295=8'd0;img296=8'd8;img297=8'd26;img298=8'd3;img299=8'd14;img300=8'd101;img301=8'd127;img302=8'd127;img303=8'd78;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd40;img314=8'd127;img315=8'd127;img316=8'd127;img317=8'd127;img318=8'd127;img319=8'd127;img320=8'd105;img321=8'd21;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd18;img329=8'd127;img330=8'd127;img331=8'd98;img332=8'd17;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd43;img342=8'd127;img343=8'd127;img344=8'd127;img345=8'd127;img346=8'd127;img347=8'd117;img348=8'd21;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd21;img357=8'd127;img358=8'd127;img359=8'd127;img360=8'd39;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd127;img370=8'd127;img371=8'd127;img372=8'd127;img373=8'd127;img374=8'd127;img375=8'd83;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd106;img385=8'd127;img386=8'd127;img387=8'd127;img388=8'd39;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd127;img398=8'd127;img399=8'd127;img400=8'd127;img401=8'd127;img402=8'd86;img403=8'd9;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd106;img413=8'd127;img414=8'd127;img415=8'd127;img416=8'd39;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd127;img426=8'd127;img427=8'd127;img428=8'd127;img429=8'd105;img430=8'd2;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd21;img438=8'd115;img439=8'd123;img440=8'd126;img441=8'd127;img442=8'd127;img443=8'd80;img444=8'd2;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd127;img454=8'd127;img455=8'd127;img456=8'd127;img457=8'd105;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd50;img464=8'd75;img465=8'd105;img466=8'd127;img467=8'd127;img468=8'd127;img469=8'd127;img470=8'd121;img471=8'd33;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd128;img482=8'd127;img483=8'd127;img484=8'd127;img485=8'd109;img486=8'd27;img487=8'd27;img488=8'd27;img489=8'd90;img490=8'd114;img491=8'd122;img492=8'd127;img493=8'd127;img494=8'd127;img495=8'd127;img496=8'd127;img497=8'd127;img498=8'd39;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd82;img510=8'd127;img511=8'd127;img512=8'd127;img513=8'd127;img514=8'd127;img515=8'd127;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd127;img520=8'd127;img521=8'd127;img522=8'd127;img523=8'd127;img524=8'd127;img525=8'd97;img526=8'd15;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd40;img538=8'd127;img539=8'd127;img540=8'd127;img541=8'd127;img542=8'd127;img543=8'd127;img544=8'd127;img545=8'd127;img546=8'd127;img547=8'd127;img548=8'd127;img549=8'd127;img550=8'd127;img551=8'd117;img552=8'd97;img553=8'd12;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd22;img566=8'd105;img567=8'd127;img568=8'd127;img569=8'd127;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd115;img579=8'd34;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd19;img595=8'd114;img596=8'd127;img597=8'd127;img598=8'd127;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd124;img605=8'd118;img606=8'd33;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd20;img624=8'd105;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd127;img629=8'd127;img630=8'd127;img631=8'd95;img632=8'd57;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd22;img653=8'd54;img654=8'd127;img655=8'd127;img656=8'd90;img657=8'd39;img658=8'd39;img659=8'd14;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd11;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd6;img235=8'd46;img236=8'd87;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd31;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd71;img259=8'd0;img260=8'd11;img261=8'd51;img262=8'd107;img263=8'd126;img264=8'd117;img265=8'd76;img266=8'd66;img267=8'd66;img268=8'd127;img269=8'd126;img270=8'd71;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd82;img286=8'd76;img287=8'd76;img288=8'd107;img289=8'd117;img290=8'd92;img291=8'd51;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd66;img297=8'd127;img298=8'd128;img299=8'd25;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd41;img313=8'd122;img314=8'd127;img315=8'd126;img316=8'd66;img317=8'd15;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd5;img325=8'd106;img326=8'd127;img327=8'd66;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd62;img341=8'd102;img342=8'd51;img343=8'd10;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd102;img354=8'd128;img355=8'd76;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd81;img382=8'd127;img383=8'd76;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd51;img410=8'd127;img411=8'd76;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd51;img438=8'd127;img439=8'd76;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd82;img466=8'd127;img467=8'd46;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd102;img494=8'd127;img495=8'd25;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd102;img522=8'd102;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd11;img549=8'd112;img550=8'd61;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd36;img577=8'd127;img578=8'd51;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd117;img605=8'd126;img606=8'd51;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd127;img633=8'd117;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd21;img660=8'd127;img661=8'd76;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd62;img688=8'd127;img689=8'd25;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd11;img715=8'd112;img716=8'd117;img717=8'd15;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd26;img743=8'd127;img744=8'd92;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd26;img771=8'd126;img772=8'd10;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd111;img153=8'd58;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd26;img180=8'd127;img181=8'd74;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd11;img187=8'd115;img188=8'd67;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd84;img208=8'd127;img209=8'd58;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd12;img215=8'd127;img216=8'd92;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd26;img235=8'd117;img236=8'd127;img237=8'd41;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd46;img243=8'd127;img244=8'd92;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd7;img262=8'd111;img263=8'd127;img264=8'd80;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd71;img271=8'd127;img272=8'd64;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd57;img290=8'd127;img291=8'd127;img292=8'd38;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd104;img299=8'd127;img300=8'd47;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd8;img317=8'd116;img318=8'd127;img319=8'd51;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd104;img327=8'd127;img328=8'd9;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd115;img345=8'd127;img346=8'd101;img347=8'd10;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd17;img354=8'd120;img355=8'd127;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd4;img371=8'd85;img372=8'd127;img373=8'd127;img374=8'd23;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd24;img382=8'd127;img383=8'd127;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd12;img399=8'd127;img400=8'd127;img401=8'd127;img402=8'd117;img403=8'd82;img404=8'd24;img405=8'd24;img406=8'd13;img407=8'd0;img408=8'd0;img409=8'd65;img410=8'd127;img411=8'd127;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd11;img427=8'd123;img428=8'd127;img429=8'd127;img430=8'd127;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd116;img435=8'd87;img436=8'd104;img437=8'd116;img438=8'd127;img439=8'd89;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd42;img456=8'd81;img457=8'd106;img458=8'd110;img459=8'd110;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd127;img466=8'd122;img467=8'd35;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd47;img489=8'd71;img490=8'd71;img491=8'd47;img492=8'd85;img493=8'd127;img494=8'd115;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd77;img521=8'd127;img522=8'd107;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd85;img549=8'd127;img550=8'd69;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd110;img577=8'd127;img578=8'd69;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd30;img604=8'd128;img605=8'd127;img606=8'd40;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd47;img632=8'd127;img633=8'd127;img634=8'd23;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd26;img660=8'd127;img661=8'd108;img662=8'd5;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd93;img689=8'd53;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd16;img150=8'd128;img151=8'd127;img152=8'd128;img153=8'd127;img154=8'd127;img155=8'd127;img156=8'd79;img157=8'd65;img158=8'd44;img159=8'd1;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd16;img178=8'd127;img179=8'd127;img180=8'd127;img181=8'd127;img182=8'd127;img183=8'd127;img184=8'd127;img185=8'd127;img186=8'd127;img187=8'd54;img188=8'd1;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd7;img206=8'd65;img207=8'd119;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd127;img216=8'd15;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd28;img236=8'd127;img237=8'd124;img238=8'd84;img239=8'd118;img240=8'd127;img241=8'd127;img242=8'd127;img243=8'd127;img244=8'd52;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd3;img263=8'd89;img264=8'd127;img265=8'd91;img266=8'd0;img267=8'd14;img268=8'd67;img269=8'd124;img270=8'd127;img271=8'd127;img272=8'd108;img273=8'd8;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd3;img290=8'd65;img291=8'd127;img292=8'd111;img293=8'd14;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd93;img298=8'd127;img299=8'd127;img300=8'd127;img301=8'd12;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd16;img318=8'd127;img319=8'd127;img320=8'd61;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd34;img326=8'd123;img327=8'd127;img328=8'd127;img329=8'd53;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd59;img346=8'd127;img347=8'd100;img348=8'd13;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd94;img355=8'd127;img356=8'd127;img357=8'd74;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd23;img373=8'd113;img374=8'd123;img375=8'd34;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd44;img383=8'd127;img384=8'd127;img385=8'd74;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd75;img401=8'd127;img402=8'd93;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd44;img411=8'd127;img412=8'd127;img413=8'd74;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd8;img428=8'd114;img429=8'd127;img430=8'd47;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd44;img439=8'd127;img440=8'd127;img441=8'd74;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd10;img456=8'd127;img457=8'd127;img458=8'd47;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd44;img467=8'd127;img468=8'd127;img469=8'd74;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd10;img484=8'd127;img485=8'd127;img486=8'd47;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd44;img495=8'd127;img496=8'd127;img497=8'd55;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd10;img512=8'd127;img513=8'd127;img514=8'd67;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd44;img523=8'd127;img524=8'd110;img525=8'd8;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd10;img540=8'd127;img541=8'd127;img542=8'd115;img543=8'd16;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd66;img551=8'd127;img552=8'd77;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd10;img568=8'd127;img569=8'd127;img570=8'd127;img571=8'd117;img572=8'd60;img573=8'd0;img574=8'd37;img575=8'd50;img576=8'd50;img577=8'd100;img578=8'd124;img579=8'd109;img580=8'd17;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd1;img596=8'd80;img597=8'd127;img598=8'd127;img599=8'd127;img600=8'd125;img601=8'd115;img602=8'd124;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd127;img607=8'd55;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd48;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd127;img629=8'd127;img630=8'd127;img631=8'd127;img632=8'd127;img633=8'd127;img634=8'd59;img635=8'd2;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd1;img653=8'd21;img654=8'd127;img655=8'd127;img656=8'd127;img657=8'd127;img658=8'd127;img659=8'd127;img660=8'd127;img661=8'd60;img662=8'd1;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd8;img682=8'd26;img683=8'd44;img684=8'd107;img685=8'd83;img686=8'd50;img687=8'd3;img688=8'd3;img689=8'd1;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd109;img124=8'd127;img125=8'd6;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd109;img152=8'd126;img153=8'd46;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd100;img180=8'd126;img181=8'd126;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd40;img208=8'd102;img209=8'd125;img210=8'd12;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd40;img237=8'd125;img238=8'd75;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd55;img265=8'd126;img266=8'd121;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd104;img293=8'd126;img294=8'd121;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd63;img321=8'd126;img322=8'd121;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd80;img349=8'd126;img350=8'd121;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd115;img377=8'd126;img378=8'd127;img379=8'd52;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd27;img405=8'd92;img406=8'd128;img407=8'd86;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd61;img434=8'd127;img435=8'd114;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd61;img462=8'd127;img463=8'd114;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd61;img490=8'd127;img491=8'd114;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd61;img518=8'd127;img519=8'd114;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd107;img546=8'd127;img547=8'd118;img548=8'd14;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd101;img574=8'd127;img575=8'd126;img576=8'd48;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd61;img602=8'd127;img603=8'd126;img604=8'd48;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd61;img630=8'd127;img631=8'd126;img632=8'd48;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd32;img658=8'd98;img659=8'd121;img660=8'd25;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd11;img176=8'd57;img177=8'd97;img178=8'd127;img179=8'd127;img180=8'd127;img181=8'd127;img182=8'd127;img183=8'd86;img184=8'd41;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd92;img204=8'd127;img205=8'd126;img206=8'd127;img207=8'd126;img208=8'd127;img209=8'd126;img210=8'd127;img211=8'd126;img212=8'd122;img213=8'd20;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd102;img232=8'd128;img233=8'd117;img234=8'd92;img235=8'd51;img236=8'd102;img237=8'd102;img238=8'd117;img239=8'd127;img240=8'd127;img241=8'd76;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd41;img260=8'd76;img261=8'd25;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd21;img266=8'd97;img267=8'd126;img268=8'd127;img269=8'd56;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd6;img293=8'd107;img294=8'd127;img295=8'd127;img296=8'd102;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd62;img320=8'd107;img321=8'd126;img322=8'd127;img323=8'd126;img324=8'd41;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd26;img347=8'd127;img348=8'd127;img349=8'd127;img350=8'd127;img351=8'd76;img352=8'd11;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd5;img375=8'd106;img376=8'd127;img377=8'd126;img378=8'd127;img379=8'd116;img380=8'd112;img381=8'd61;img382=8'd41;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd62;img405=8'd112;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd36;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd10;img434=8'd25;img435=8'd66;img436=8'd107;img437=8'd126;img438=8'd127;img439=8'd96;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd11;img465=8'd81;img466=8'd127;img467=8'd127;img468=8'd51;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd11;img493=8'd102;img494=8'd127;img495=8'd126;img496=8'd31;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd66;img521=8'd127;img522=8'd127;img523=8'd46;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd11;img547=8'd71;img548=8'd127;img549=8'd126;img550=8'd117;img551=8'd15;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd21;img574=8'd107;img575=8'd127;img576=8'd127;img577=8'd107;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd82;img601=8'd122;img602=8'd127;img603=8'd126;img604=8'd86;img605=8'd5;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd6;img625=8'd87;img626=8'd87;img627=8'd127;img628=8'd128;img629=8'd127;img630=8'd112;img631=8'd41;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd66;img653=8'd126;img654=8'd127;img655=8'd126;img656=8'd127;img657=8'd86;img658=8'd10;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd77;img681=8'd127;img682=8'd122;img683=8'd102;img684=8'd41;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd46;img709=8'd96;img710=8'd61;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd102;img153=8'd97;img154=8'd15;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd102;img181=8'd127;img182=8'd66;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd51;img209=8'd127;img210=8'd76;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd51;img237=8'd127;img238=8'd76;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd21;img265=8'd127;img266=8'd127;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd127;img294=8'd126;img295=8'd41;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd76;img322=8'd127;img323=8'd102;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd76;img350=8'd126;img351=8'd102;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd46;img378=8'd127;img379=8'd107;img380=8'd5;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd5;img406=8'd106;img407=8'd127;img408=8'd25;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd102;img435=8'd127;img436=8'd56;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd81;img463=8'd127;img464=8'd76;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd51;img491=8'd127;img492=8'd76;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd51;img519=8'd127;img520=8'd96;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd51;img547=8'd127;img548=8'd127;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd51;img575=8'd127;img576=8'd126;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd21;img603=8'd128;img604=8'd127;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd127;img632=8'd126;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd87;img660=8'd127;img661=8'd31;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd26;img688=8'd126;img689=8'd51;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd50;img149=8'd127;img150=8'd127;img151=8'd127;img152=8'd127;img153=8'd109;img154=8'd59;img155=8'd21;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd89;img176=8'd124;img177=8'd127;img178=8'd127;img179=8'd127;img180=8'd127;img181=8'd127;img182=8'd127;img183=8'd70;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd32;img203=8'd122;img204=8'd127;img205=8'd104;img206=8'd89;img207=8'd89;img208=8'd28;img209=8'd50;img210=8'd127;img211=8'd125;img212=8'd46;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd10;img231=8'd83;img232=8'd90;img233=8'd13;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd35;img238=8'd127;img239=8'd127;img240=8'd55;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd35;img266=8'd127;img267=8'd125;img268=8'd48;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd7;img293=8'd77;img294=8'd127;img295=8'd72;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd29;img320=8'd120;img321=8'd127;img322=8'd127;img323=8'd45;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd3;img346=8'd56;img347=8'd124;img348=8'd127;img349=8'd127;img350=8'd114;img351=8'd21;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd16;img373=8'd114;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd111;img380=8'd44;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd18;img401=8'd127;img402=8'd127;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd126;img409=8'd103;img410=8'd24;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd14;img429=8'd103;img430=8'd103;img431=8'd103;img432=8'd41;img433=8'd34;img434=8'd34;img435=8'd94;img436=8'd127;img437=8'd127;img438=8'd113;img439=8'd26;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd29;img464=8'd84;img465=8'd127;img466=8'd127;img467=8'd112;img468=8'd18;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd2;img493=8'd88;img494=8'd127;img495=8'd127;img496=8'd29;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd87;img523=8'd127;img524=8'd111;img525=8'd19;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd52;img551=8'd127;img552=8'd127;img553=8'd38;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd21;img578=8'd114;img579=8'd127;img580=8'd127;img581=8'd38;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd6;img603=8'd32;img604=8'd70;img605=8'd113;img606=8'd127;img607=8'd127;img608=8'd119;img609=8'd29;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd21;img628=8'd21;img629=8'd77;img630=8'd97;img631=8'd127;img632=8'd127;img633=8'd127;img634=8'd127;img635=8'd109;img636=8'd43;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd2;img653=8'd15;img654=8'd79;img655=8'd126;img656=8'd127;img657=8'd127;img658=8'd127;img659=8'd127;img660=8'd127;img661=8'd116;img662=8'd51;img663=8'd7;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd8;img681=8'd58;img682=8'd93;img683=8'd127;img684=8'd127;img685=8'd127;img686=8'd114;img687=8'd58;img688=8'd57;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd8;img123=8'd1;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd94;img151=8'd88;img152=8'd38;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd11;img164=8'd2;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd69;img179=8'd127;img180=8'd57;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd67;img192=8'd70;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd54;img207=8'd127;img208=8'd57;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd35;img219=8'd124;img220=8'd127;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd107;img235=8'd127;img236=8'd57;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd67;img247=8'd127;img248=8'd102;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd22;img262=8'd120;img263=8'd127;img264=8'd57;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd101;img275=8'd127;img276=8'd39;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd51;img290=8'd127;img291=8'd127;img292=8'd51;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd4;img302=8'd104;img303=8'd123;img304=8'd8;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd6;img317=8'd108;img318=8'd127;img319=8'd87;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd43;img330=8'd127;img331=8'd77;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd78;img345=8'd127;img346=8'd127;img347=8'd24;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd92;img358=8'd127;img359=8'd77;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd39;img372=8'd120;img373=8'd127;img374=8'd111;img375=8'd4;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd8;img385=8'd103;img386=8'd127;img387=8'd77;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd7;img399=8'd102;img400=8'd127;img401=8'd127;img402=8'd24;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd24;img413=8'd127;img414=8'd127;img415=8'd27;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd18;img427=8'd127;img428=8'd127;img429=8'd87;img430=8'd2;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd24;img441=8'd127;img442=8'd127;img443=8'd18;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd36;img454=8'd102;img455=8'd127;img456=8'd109;img457=8'd13;img458=8'd0;img459=8'd1;img460=8'd6;img461=8'd6;img462=8'd6;img463=8'd4;img464=8'd6;img465=8'd6;img466=8'd1;img467=8'd0;img468=8'd24;img469=8'd127;img470=8'd87;img471=8'd1;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd75;img482=8'd127;img483=8'd127;img484=8'd113;img485=8'd74;img486=8'd74;img487=8'd76;img488=8'd127;img489=8'd127;img490=8'd128;img491=8'd103;img492=8'd127;img493=8'd127;img494=8'd45;img495=8'd7;img496=8'd59;img497=8'd127;img498=8'd79;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd117;img510=8'd127;img511=8'd127;img512=8'd127;img513=8'd127;img514=8'd127;img515=8'd127;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd109;img520=8'd113;img521=8'd106;img522=8'd127;img523=8'd102;img524=8'd112;img525=8'd127;img526=8'd27;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd54;img538=8'd127;img539=8'd127;img540=8'd112;img541=8'd101;img542=8'd95;img543=8'd95;img544=8'd62;img545=8'd36;img546=8'd36;img547=8'd9;img548=8'd14;img549=8'd4;img550=8'd35;img551=8'd89;img552=8'd127;img553=8'd104;img554=8'd8;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd2;img566=8'd27;img567=8'd27;img568=8'd14;img569=8'd5;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd74;img580=8'd127;img581=8'd75;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd11;img608=8'd18;img609=8'd5;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd114;img176=8'd106;img177=8'd45;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd26;img185=8'd61;img186=8'd61;img187=8'd113;img188=8'd127;img189=8'd116;img190=8'd22;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd31;img204=8'd118;img205=8'd125;img206=8'd120;img207=8'd120;img208=8'd120;img209=8'd120;img210=8'd120;img211=8'd121;img212=8'd123;img213=8'd126;img214=8'd126;img215=8'd126;img216=8'd126;img217=8'd126;img218=8'd47;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd32;img233=8'd92;img234=8'd126;img235=8'd126;img236=8'd126;img237=8'd126;img238=8'd126;img239=8'd127;img240=8'd126;img241=8'd126;img242=8'd126;img243=8'd126;img244=8'd126;img245=8'd126;img246=8'd47;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd6;img262=8'd20;img263=8'd20;img264=8'd27;img265=8'd48;img266=8'd20;img267=8'd20;img268=8'd20;img269=8'd20;img270=8'd110;img271=8'd126;img272=8'd126;img273=8'd99;img274=8'd32;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd38;img298=8'd122;img299=8'd126;img300=8'd105;img301=8'd9;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd61;img326=8'd126;img327=8'd126;img328=8'd99;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd48;img353=8'd122;img354=8'd126;img355=8'd126;img356=8'd89;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd7;img380=8'd121;img381=8'd126;img382=8'd126;img383=8'd63;img384=8'd12;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd4;img407=8'd99;img408=8'd126;img409=8'd126;img410=8'd124;img411=8'd25;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd4;img434=8'd98;img435=8'd127;img436=8'd126;img437=8'd126;img438=8'd51;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd7;img461=8'd99;img462=8'd127;img463=8'd128;img464=8'd127;img465=8'd80;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd9;img488=8'd62;img489=8'd126;img490=8'd126;img491=8'd127;img492=8'd126;img493=8'd52;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd45;img516=8'd126;img517=8'd126;img518=8'd126;img519=8'd127;img520=8'd19;img521=8'd2;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd9;img543=8'd99;img544=8'd126;img545=8'd126;img546=8'd105;img547=8'd55;img548=8'd1;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd9;img570=8'd88;img571=8'd126;img572=8'd126;img573=8'd124;img574=8'd44;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd9;img597=8'd54;img598=8'd126;img599=8'd126;img600=8'd126;img601=8'd70;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd86;img625=8'd126;img626=8'd126;img627=8'd126;img628=8'd117;img629=8'd17;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd5;img652=8'd109;img653=8'd126;img654=8'd126;img655=8'd126;img656=8'd70;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd45;img680=8'd125;img681=8'd126;img682=8'd126;img683=8'd111;img684=8'd20;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd107;img709=8'd109;img710=8'd109;img711=8'd40;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd18;img125=8'd63;img126=8'd96;img127=8'd109;img128=8'd128;img129=8'd127;img130=8'd127;img131=8'd121;img132=8'd26;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd102;img152=8'd125;img153=8'd127;img154=8'd127;img155=8'd127;img156=8'd127;img157=8'd127;img158=8'd127;img159=8'd127;img160=8'd125;img161=8'd118;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd44;img178=8'd121;img179=8'd126;img180=8'd127;img181=8'd113;img182=8'd71;img183=8'd25;img184=8'd6;img185=8'd6;img186=8'd6;img187=8'd53;img188=8'd127;img189=8'd127;img190=8'd56;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd48;img205=8'd113;img206=8'd127;img207=8'd84;img208=8'd57;img209=8'd7;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd8;img216=8'd106;img217=8'd127;img218=8'd59;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd46;img232=8'd119;img233=8'd127;img234=8'd85;img235=8'd14;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd75;img245=8'd127;img246=8'd59;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd49;img259=8'd126;img260=8'd109;img261=8'd24;img262=8'd3;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd75;img273=8'd127;img274=8'd59;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd56;img287=8'd127;img288=8'd56;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd5;img300=8'd92;img301=8'd121;img302=8'd9;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd10;img315=8'd23;img316=8'd3;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd34;img328=8'd127;img329=8'd120;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd14;img355=8'd117;img356=8'd124;img357=8'd53;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd22;img382=8'd79;img383=8'd127;img384=8'd66;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd6;img409=8'd95;img410=8'd127;img411=8'd102;img412=8'd14;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd6;img436=8'd78;img437=8'd127;img438=8'd123;img439=8'd39;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd6;img463=8'd78;img464=8'd127;img465=8'd101;img466=8'd34;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd6;img490=8'd78;img491=8'd127;img492=8'd113;img493=8'd36;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd15;img513=8'd17;img514=8'd17;img515=8'd70;img516=8'd82;img517=8'd93;img518=8'd127;img519=8'd113;img520=8'd19;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd6;img539=8'd41;img540=8'd122;img541=8'd127;img542=8'd127;img543=8'd127;img544=8'd127;img545=8'd127;img546=8'd127;img547=8'd127;img548=8'd93;img549=8'd35;img550=8'd12;img551=8'd0;img552=8'd0;img553=8'd11;img554=8'd78;img555=8'd39;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd40;img566=8'd98;img567=8'd127;img568=8'd127;img569=8'd127;img570=8'd127;img571=8'd127;img572=8'd124;img573=8'd117;img574=8'd83;img575=8'd124;img576=8'd127;img577=8'd127;img578=8'd120;img579=8'd75;img580=8'd37;img581=8'd72;img582=8'd52;img583=8'd26;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd4;img593=8'd124;img594=8'd127;img595=8'd127;img596=8'd127;img597=8'd127;img598=8'd127;img599=8'd121;img600=8'd53;img601=8'd0;img602=8'd0;img603=8'd54;img604=8'd121;img605=8'd127;img606=8'd127;img607=8'd127;img608=8'd123;img609=8'd80;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd29;img621=8'd125;img622=8'd127;img623=8'd127;img624=8'd127;img625=8'd124;img626=8'd68;img627=8'd11;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd11;img633=8'd59;img634=8'd92;img635=8'd92;img636=8'd24;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd61;img650=8'd62;img651=8'd88;img652=8'd68;img653=8'd8;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd31;img203=8'd78;img204=8'd74;img205=8'd45;img206=8'd41;img207=8'd78;img208=8'd128;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd108;img213=8'd78;img214=8'd74;img215=8'd21;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd13;img230=8'd104;img231=8'd127;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd123;img236=8'd117;img237=8'd98;img238=8'd117;img239=8'd117;img240=8'd117;img241=8'd123;img242=8'd127;img243=8'd121;img244=8'd12;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd83;img258=8'd127;img259=8'd127;img260=8'd127;img261=8'd127;img262=8'd64;img263=8'd24;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd24;img270=8'd113;img271=8'd127;img272=8'd44;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd2;img284=8'd87;img285=8'd126;img286=8'd127;img287=8'd122;img288=8'd62;img289=8'd10;img290=8'd1;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd107;img299=8'd127;img300=8'd10;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd66;img312=8'd127;img313=8'd127;img314=8'd89;img315=8'd23;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd23;img326=8'd122;img327=8'd127;img328=8'd10;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd64;img340=8'd98;img341=8'd45;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd90;img354=8'd127;img355=8'd76;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd4;img381=8'd127;img382=8'd126;img383=8'd36;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd83;img409=8'd127;img410=8'd83;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd19;img436=8'd124;img437=8'd127;img438=8'd23;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd39;img464=8'd127;img465=8'd86;img466=8'd5;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd10;img491=8'd120;img492=8'd127;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd1;img518=8'd46;img519=8'd127;img520=8'd127;img521=8'd108;img522=8'd107;img523=8'd107;img524=8'd91;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd10;img545=8'd84;img546=8'd127;img547=8'd127;img548=8'd127;img549=8'd127;img550=8'd127;img551=8'd127;img552=8'd107;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd101;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd93;img577=8'd59;img578=8'd17;img579=8'd10;img580=8'd8;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd60;img601=8'd37;img602=8'd97;img603=8'd119;img604=8'd18;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd40;img630=8'd127;img631=8'd107;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd59;img658=8'd127;img659=8'd84;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd59;img686=8'd127;img687=8'd59;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd59;img714=8'd127;img715=8'd59;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd36;img742=8'd97;img743=8'd17;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd7;img152=8'd109;img153=8'd105;img154=8'd31;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd3;img180=8'd95;img181=8'd126;img182=8'd93;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd85;img209=8'd126;img210=8'd108;img211=8'd3;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd85;img237=8'd126;img238=8'd127;img239=8'd32;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd85;img265=8'd126;img266=8'd127;img267=8'd32;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd55;img293=8'd127;img294=8'd127;img295=8'd84;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd32;img321=8'd126;img322=8'd127;img323=8'd84;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd30;img349=8'd125;img350=8'd127;img351=8'd105;img352=8'd6;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd106;img378=8'd127;img379=8'd126;img380=8'd11;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd106;img406=8'd127;img407=8'd126;img408=8'd11;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd106;img434=8'd128;img435=8'd127;img436=8'd11;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd106;img462=8'd127;img463=8'd126;img464=8'd11;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd106;img490=8'd127;img491=8'd126;img492=8'd11;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd84;img518=8'd127;img519=8'd126;img520=8'd11;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd106;img546=8'd127;img547=8'd126;img548=8'd11;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd106;img574=8'd128;img575=8'd127;img576=8'd11;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd66;img602=8'd127;img603=8'd126;img604=8'd11;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd53;img630=8'd127;img631=8'd126;img632=8'd11;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd53;img658=8'd127;img659=8'd126;img660=8'd11;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd9;img686=8'd105;img687=8'd91;img688=8'd2;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd25;img126=8'd85;img127=8'd127;img128=8'd30;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd18;img152=8'd96;img153=8'd123;img154=8'd127;img155=8'd127;img156=8'd88;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd2;img178=8'd35;img179=8'd121;img180=8'd127;img181=8'd118;img182=8'd117;img183=8'd127;img184=8'd91;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd12;img205=8'd92;img206=8'd127;img207=8'd122;img208=8'd50;img209=8'd14;img210=8'd55;img211=8'd127;img212=8'd91;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd10;img232=8'd103;img233=8'd124;img234=8'd49;img235=8'd13;img236=8'd0;img237=8'd0;img238=8'd55;img239=8'd127;img240=8'd75;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd20;img260=8'd52;img261=8'd10;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd55;img267=8'd127;img268=8'd17;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd55;img295=8'd117;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd16;img322=8'd107;img323=8'd75;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd67;img350=8'd100;img351=8'd8;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd10;img377=8'd116;img378=8'd72;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd73;img405=8'd122;img406=8'd36;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd8;img432=8'd101;img433=8'd66;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd82;img460=8'd113;img461=8'd16;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd6;img470=8'd61;img471=8'd103;img472=8'd24;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd40;img487=8'd128;img488=8'd64;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd8;img496=8'd42;img497=8'd108;img498=8'd125;img499=8'd72;img500=8'd6;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd4;img514=8'd104;img515=8'd114;img516=8'd19;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd10;img522=8'd68;img523=8'd119;img524=8'd127;img525=8'd114;img526=8'd32;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd68;img542=8'd127;img543=8'd33;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd27;img548=8'd95;img549=8'd127;img550=8'd127;img551=8'd99;img552=8'd59;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd11;img569=8'd116;img570=8'd91;img571=8'd0;img572=8'd16;img573=8'd51;img574=8'd92;img575=8'd125;img576=8'd120;img577=8'd90;img578=8'd48;img579=8'd2;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd64;img597=8'd127;img598=8'd50;img599=8'd64;img600=8'd116;img601=8'd127;img602=8'd126;img603=8'd93;img604=8'd30;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd2;img624=8'd111;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd127;img629=8'd96;img630=8'd35;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd28;img652=8'd127;img653=8'd127;img654=8'd94;img655=8'd53;img656=8'd36;img657=8'd6;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd33;img127=8'd111;img128=8'd15;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd16;img154=8'd112;img155=8'd127;img156=8'd64;img157=8'd5;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd33;img182=8'd127;img183=8'd127;img184=8'd127;img185=8'd87;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd91;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd87;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd91;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd79;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd91;img266=8'd127;img267=8'd127;img268=8'd122;img269=8'd21;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd17;img293=8'd115;img294=8'd127;img295=8'd127;img296=8'd90;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd68;img321=8'd127;img322=8'd127;img323=8'd127;img324=8'd78;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd5;img348=8'd96;img349=8'd127;img350=8'd127;img351=8'd127;img352=8'd28;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd22;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd28;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd22;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd118;img408=8'd21;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd22;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd93;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd22;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd43;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd22;img488=8'd127;img489=8'd127;img490=8'd101;img491=8'd6;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd12;img516=8'd108;img517=8'd127;img518=8'd123;img519=8'd50;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd14;img544=8'd112;img545=8'd127;img546=8'd127;img547=8'd93;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd10;img572=8'd104;img573=8'd127;img574=8'd127;img575=8'd93;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd12;img600=8'd108;img601=8'd127;img602=8'd127;img603=8'd93;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd12;img628=8'd109;img629=8'd127;img630=8'd127;img631=8'd93;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd57;img657=8'd128;img658=8'd128;img659=8'd63;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd81;img126=8'd16;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd109;img154=8'd76;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd67;img182=8'd116;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd39;img210=8'd116;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd33;img238=8'd117;img239=8'd5;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd127;img267=8'd27;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd127;img295=8'd27;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd127;img323=8'd27;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd127;img351=8'd47;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd127;img379=8'd42;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd16;img406=8'd128;img407=8'd39;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd39;img434=8'd127;img435=8'd27;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd39;img462=8'd117;img463=8'd4;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd64;img490=8'd116;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd83;img518=8'd116;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd116;img546=8'd106;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd116;img574=8'd76;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd4;img601=8'd117;img602=8'd39;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd27;img629=8'd127;img630=8'd19;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd51;img657=8'd127;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd11;img208=8'd49;img209=8'd91;img210=8'd127;img211=8'd128;img212=8'd111;img213=8'd53;img214=8'd2;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd14;img233=8'd64;img234=8'd107;img235=8'd123;img236=8'd127;img237=8'd127;img238=8'd123;img239=8'd120;img240=8'd127;img241=8'd127;img242=8'd47;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd14;img259=8'd76;img260=8'd120;img261=8'd127;img262=8'd127;img263=8'd111;img264=8'd102;img265=8'd95;img266=8'd35;img267=8'd14;img268=8'd108;img269=8'd127;img270=8'd49;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd22;img287=8'd124;img288=8'd127;img289=8'd117;img290=8'd20;img291=8'd8;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd48;img297=8'd127;img298=8'd56;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd61;img316=8'd36;img317=8'd17;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd38;img325=8'd127;img326=8'd94;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd47;img353=8'd127;img354=8'd75;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd62;img381=8'd127;img382=8'd20;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd3;img408=8'd102;img409=8'd87;img410=8'd1;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd51;img436=8'd127;img437=8'd61;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd20;img462=8'd112;img463=8'd103;img464=8'd127;img465=8'd58;img466=8'd17;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd20;img490=8'd124;img491=8'd127;img492=8'd127;img493=8'd127;img494=8'd121;img495=8'd96;img496=8'd36;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd70;img519=8'd127;img520=8'd127;img521=8'd124;img522=8'd105;img523=8'd127;img524=8'd107;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd2;img546=8'd93;img547=8'd104;img548=8'd36;img549=8'd25;img550=8'd37;img551=8'd96;img552=8'd67;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd67;img574=8'd127;img575=8'd60;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd8;img601=8'd99;img602=8'd84;img603=8'd1;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd70;img629=8'd113;img630=8'd22;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd26;img656=8'd117;img657=8'd53;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd81;img684=8'd114;img685=8'd9;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd114;img712=8'd62;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd84;img740=8'd3;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd61;img177=8'd128;img178=8'd83;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd35;img186=8'd127;img187=8'd90;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd66;img205=8'd127;img206=8'd77;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd53;img214=8'd127;img215=8'd125;img216=8'd25;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd108;img233=8'd127;img234=8'd53;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd70;img242=8'd127;img243=8'd120;img244=8'd19;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd7;img260=8'd113;img261=8'd127;img262=8'd42;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd43;img269=8'd117;img270=8'd127;img271=8'd108;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd29;img288=8'd127;img289=8'd127;img290=8'd23;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd4;img296=8'd93;img297=8'd127;img298=8'd127;img299=8'd103;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd29;img316=8'd127;img317=8'd127;img318=8'd5;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd73;img324=8'd127;img325=8'd127;img326=8'd127;img327=8'd60;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd75;img344=8'd127;img345=8'd127;img346=8'd5;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd64;img351=8'd126;img352=8'd127;img353=8'd127;img354=8'd120;img355=8'd11;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd77;img372=8'd127;img373=8'd127;img374=8'd5;img375=8'd0;img376=8'd0;img377=8'd46;img378=8'd123;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd91;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd53;img400=8'd121;img401=8'd127;img402=8'd20;img403=8'd0;img404=8'd14;img405=8'd122;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd75;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd81;img429=8'd127;img430=8'd85;img431=8'd50;img432=8'd122;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd127;img437=8'd126;img438=8'd35;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd34;img457=8'd88;img458=8'd127;img459=8'd127;img460=8'd127;img461=8'd123;img462=8'd84;img463=8'd127;img464=8'd127;img465=8'd101;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd50;img487=8'd89;img488=8'd73;img489=8'd18;img490=8'd55;img491=8'd127;img492=8'd127;img493=8'd74;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd103;img519=8'd127;img520=8'd127;img521=8'd66;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd65;img547=8'd127;img548=8'd110;img549=8'd6;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd87;img575=8'd127;img576=8'd105;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd78;img603=8'd127;img604=8'd62;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd93;img631=8'd127;img632=8'd58;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd103;img659=8'd127;img660=8'd58;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd97;img687=8'd127;img688=8'd58;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd14;img715=8'd96;img716=8'd58;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd21;img127=8'd51;img128=8'd51;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd41;img155=8'd107;img156=8'd127;img157=8'd82;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd16;img184=8'd116;img185=8'd112;img186=8'd10;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd102;img213=8'd122;img214=8'd20;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd21;img240=8'd122;img241=8'd81;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd36;img268=8'd127;img269=8'd21;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd21;img295=8'd117;img296=8'd106;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd6;img322=8'd87;img323=8'd112;img324=8'd10;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd66;img350=8'd126;img351=8'd81;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd11;img377=8'd127;img378=8'd96;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd11;img404=8'd102;img405=8'd117;img406=8'd25;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd66;img432=8'd127;img433=8'd51;img434=8'd0;img435=8'd16;img436=8'd26;img437=8'd26;img438=8'd26;img439=8'd57;img440=8'd56;img441=8'd57;img442=8'd76;img443=8'd66;img444=8'd5;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd41;img459=8'd127;img460=8'd126;img461=8'd112;img462=8'd102;img463=8'd117;img464=8'd126;img465=8'd127;img466=8'd126;img467=8'd127;img468=8'd126;img469=8'd127;img470=8'd126;img471=8'd127;img472=8'd46;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd6;img484=8'd26;img485=8'd87;img486=8'd127;img487=8'd127;img488=8'd127;img489=8'd127;img490=8'd107;img491=8'd51;img492=8'd51;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd82;img500=8'd102;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd62;img511=8'd107;img512=8'd126;img513=8'd127;img514=8'd126;img515=8'd96;img516=8'd56;img517=8'd25;img518=8'd5;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd20;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd87;img538=8'd127;img539=8'd128;img540=8'd127;img541=8'd112;img542=8'd20;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd127;img566=8'd126;img567=8'd127;img568=8'd65;img569=8'd10;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd51;img594=8'd51;img595=8'd21;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd12;img122=8'd76;img123=8'd128;img124=8'd127;img125=8'd82;img126=8'd16;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd12;img149=8'd106;img150=8'd127;img151=8'd127;img152=8'd127;img153=8'd127;img154=8'd34;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd78;img177=8'd121;img178=8'd76;img179=8'd68;img180=8'd124;img181=8'd127;img182=8'd93;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd70;img205=8'd42;img206=8'd0;img207=8'd0;img208=8'd81;img209=8'd124;img210=8'd96;img211=8'd3;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd4;img237=8'd97;img238=8'd127;img239=8'd28;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd28;img265=8'd127;img266=8'd127;img267=8'd28;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd39;img293=8'd127;img294=8'd104;img295=8'd10;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd90;img321=8'd127;img322=8'd93;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd18;img348=8'd116;img349=8'd127;img350=8'd100;img351=8'd28;img352=8'd6;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd25;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd80;img381=8'd21;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd19;img404=8'd93;img405=8'd118;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd95;img410=8'd5;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd21;img434=8'd45;img435=8'd101;img436=8'd127;img437=8'd127;img438=8'd103;img439=8'd12;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd8;img464=8'd107;img465=8'd127;img466=8'd127;img467=8'd15;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd103;img493=8'd127;img494=8'd127;img495=8'd15;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd13;img519=8'd65;img520=8'd123;img521=8'd127;img522=8'd110;img523=8'd10;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd37;img546=8'd101;img547=8'd127;img548=8'd127;img549=8'd110;img550=8'd19;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd49;img572=8'd115;img573=8'd124;img574=8'd127;img575=8'd127;img576=8'd84;img577=8'd19;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd48;img599=8'd124;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd65;img604=8'd2;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd84;img627=8'd127;img628=8'd127;img629=8'd127;img630=8'd65;img631=8'd2;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd54;img655=8'd127;img656=8'd113;img657=8'd19;img658=8'd1;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd82;img153=8'd97;img154=8'd76;img155=8'd46;img156=8'd26;img157=8'd26;img158=8'd26;img159=8'd26;img160=8'd16;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd11;img180=8'd112;img181=8'd127;img182=8'd126;img183=8'd127;img184=8'd126;img185=8'd127;img186=8'd126;img187=8'd127;img188=8'd96;img189=8'd41;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd26;img208=8'd127;img209=8'd51;img210=8'd0;img211=8'd11;img212=8'd51;img213=8'd31;img214=8'd51;img215=8'd51;img216=8'd31;img217=8'd92;img218=8'd20;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd26;img236=8'd126;img237=8'd51;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd31;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd26;img264=8'd127;img265=8'd51;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd46;img292=8'd126;img293=8'd51;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd87;img320=8'd127;img321=8'd51;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd127;img348=8'd126;img349=8'd112;img350=8'd102;img351=8'd102;img352=8'd102;img353=8'd41;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd62;img375=8'd127;img376=8'd127;img377=8'd112;img378=8'd102;img379=8'd102;img380=8'd112;img381=8'd127;img382=8'd36;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd21;img402=8'd122;img403=8'd127;img404=8'd65;img405=8'd10;img406=8'd0;img407=8'd0;img408=8'd10;img409=8'd127;img410=8'd116;img411=8'd21;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd76;img430=8'd127;img431=8'd92;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd66;img438=8'd127;img439=8'd51;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd26;img458=8'd76;img459=8'd10;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd26;img466=8'd126;img467=8'd51;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd11;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd57;img494=8'd127;img495=8'd51;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd41;img513=8'd92;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd97;img522=8'd126;img523=8'd51;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd102;img541=8'd92;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd11;img549=8'd127;img550=8'd127;img551=8'd21;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd11;img568=8'd112;img569=8'd51;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd11;img576=8'd102;img577=8'd127;img578=8'd65;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd102;img597=8'd62;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd21;img603=8'd87;img604=8'd127;img605=8'd102;img606=8'd10;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd81;img625=8'd112;img626=8'd51;img627=8'd11;img628=8'd51;img629=8'd82;img630=8'd122;img631=8'd127;img632=8'd86;img633=8'd10;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd21;img653=8'd117;img654=8'd127;img655=8'd128;img656=8'd127;img657=8'd128;img658=8'd86;img659=8'd41;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd15;img682=8'd66;img683=8'd96;img684=8'd56;img685=8'd25;img686=8'd5;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd76;img123=8'd127;img124=8'd84;img125=8'd5;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd13;img150=8'd111;img151=8'd126;img152=8'd126;img153=8'd33;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd99;img179=8'd126;img180=8'd126;img181=8'd94;img182=8'd7;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd70;img207=8'd126;img208=8'd126;img209=8'd126;img210=8'd45;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd35;img235=8'd124;img236=8'd126;img237=8'd126;img238=8'd71;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd97;img264=8'd126;img265=8'd126;img266=8'd115;img267=8'd20;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd35;img292=8'd126;img293=8'd126;img294=8'd126;img295=8'd106;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd5;img320=8'd118;img321=8'd126;img322=8'd126;img323=8'd113;img324=8'd7;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd61;img349=8'd126;img350=8'd126;img351=8'd127;img352=8'd39;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd3;img377=8'd98;img378=8'd126;img379=8'd127;img380=8'd101;img381=8'd10;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd94;img406=8'd127;img407=8'd128;img408=8'd127;img409=8'd22;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd79;img434=8'd126;img435=8'd127;img436=8'd126;img437=8'd61;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd39;img462=8'd126;img463=8'd127;img464=8'd126;img465=8'd96;img466=8'd2;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd2;img490=8'd106;img491=8'd127;img492=8'd126;img493=8'd126;img494=8'd58;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd56;img519=8'd127;img520=8'd126;img521=8'd126;img522=8'd96;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd36;img547=8'd127;img548=8'd126;img549=8'd126;img550=8'd119;img551=8'd16;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd100;img576=8'd126;img577=8'd126;img578=8'd126;img579=8'd70;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd63;img604=8'd126;img605=8'd126;img606=8'd126;img607=8'd99;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd17;img632=8'd126;img633=8'd126;img634=8'd126;img635=8'd58;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd3;img660=8'd55;img661=8'd117;img662=8'd122;img663=8'd25;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd38;img66=8'd87;img67=8'd113;img68=8'd128;img69=8'd93;img70=8'd27;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd111;img94=8'd42;img95=8'd34;img96=8'd37;img97=8'd93;img98=8'd122;img99=8'd61;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd48;img122=8'd6;img123=8'd0;img124=8'd0;img125=8'd4;img126=8'd57;img127=8'd121;img128=8'd49;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd4;img155=8'd57;img156=8'd111;img157=8'd12;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd12;img184=8'd110;img185=8'd84;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd36;img213=8'd112;img214=8'd1;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd22;img241=8'd125;img242=8'd42;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd91;img270=8'd83;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd109;img298=8'd83;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd6;img325=8'd121;img326=8'd83;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd33;img353=8'd127;img354=8'd49;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd33;img381=8'd127;img382=8'd19;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd36;img403=8'd40;img404=8'd51;img405=8'd10;img406=8'd0;img407=8'd0;img408=8'd83;img409=8'd91;img410=8'd1;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd10;img429=8'd80;img430=8'd121;img431=8'd123;img432=8'd123;img433=8'd121;img434=8'd60;img435=8'd30;img436=8'd127;img437=8'd48;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd94;img457=8'd112;img458=8'd18;img459=8'd0;img460=8'd3;img461=8'd58;img462=8'd122;img463=8'd127;img464=8'd104;img465=8'd3;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd14;img484=8'd122;img485=8'd52;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd41;img491=8'd127;img492=8'd109;img493=8'd9;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd32;img512=8'd127;img513=8'd16;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd39;img518=8'd122;img519=8'd107;img520=8'd113;img521=8'd100;img522=8'd8;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd19;img540=8'd127;img541=8'd25;img542=8'd0;img543=8'd28;img544=8'd47;img545=8'd123;img546=8'd107;img547=8'd15;img548=8'd21;img549=8'd114;img550=8'd101;img551=8'd29;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd2;img568=8'd96;img569=8'd121;img570=8'd115;img571=8'd127;img572=8'd127;img573=8'd84;img574=8'd15;img575=8'd0;img576=8'd0;img577=8'd20;img578=8'd67;img579=8'd122;img580=8'd92;img581=8'd35;img582=8'd16;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd11;img597=8'd69;img598=8'd87;img599=8'd47;img600=8'd6;img601=8'd2;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd1;img607=8'd51;img608=8'd105;img609=8'd120;img610=8'd27;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd2;img178=8'd56;img179=8'd67;img180=8'd41;img181=8'd1;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd2;img186=8'd50;img187=8'd84;img188=8'd107;img189=8'd10;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd43;img206=8'd127;img207=8'd127;img208=8'd127;img209=8'd6;img210=8'd0;img211=8'd0;img212=8'd2;img213=8'd64;img214=8'd127;img215=8'd127;img216=8'd127;img217=8'd18;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd28;img233=8'd116;img234=8'd127;img235=8'd127;img236=8'd119;img237=8'd5;img238=8'd0;img239=8'd0;img240=8'd19;img241=8'd127;img242=8'd127;img243=8'd127;img244=8'd127;img245=8'd56;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd91;img261=8'd127;img262=8'd127;img263=8'd127;img264=8'd72;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd19;img269=8'd127;img270=8'd127;img271=8'd127;img272=8'd127;img273=8'd67;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd32;img288=8'd117;img289=8'd127;img290=8'd127;img291=8'd127;img292=8'd29;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd19;img297=8'd127;img298=8'd127;img299=8'd127;img300=8'd127;img301=8'd18;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd6;img315=8'd97;img316=8'd127;img317=8'd127;img318=8'd127;img319=8'd127;img320=8'd12;img321=8'd0;img322=8'd2;img323=8'd43;img324=8'd101;img325=8'd127;img326=8'd127;img327=8'd127;img328=8'd127;img329=8'd18;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd19;img343=8'd127;img344=8'd127;img345=8'd127;img346=8'd127;img347=8'd127;img348=8'd51;img349=8'd43;img350=8'd105;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd127;img355=8'd127;img356=8'd92;img357=8'd4;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd71;img371=8'd127;img372=8'd127;img373=8'd127;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd127;img383=8'd127;img384=8'd33;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd53;img399=8'd127;img400=8'd127;img401=8'd127;img402=8'd127;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd94;img412=8'd3;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd19;img427=8'd127;img428=8'd127;img429=8'd127;img430=8'd127;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd90;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd18;img455=8'd124;img456=8'd121;img457=8'd75;img458=8'd110;img459=8'd121;img460=8'd121;img461=8'd121;img462=8'd122;img463=8'd127;img464=8'd127;img465=8'd128;img466=8'd127;img467=8'd88;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd26;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd3;img491=8'd96;img492=8'd127;img493=8'd127;img494=8'd127;img495=8'd30;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd73;img520=8'd127;img521=8'd127;img522=8'd127;img523=8'd39;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd5;img547=8'd109;img548=8'd127;img549=8'd127;img550=8'd127;img551=8'd90;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd21;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd127;img579=8'd76;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd113;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd127;img607=8'd30;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd50;img630=8'd127;img631=8'd127;img632=8'd127;img633=8'd127;img634=8'd127;img635=8'd30;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd61;img658=8'd127;img659=8'd127;img660=8'd127;img661=8'd127;img662=8'd115;img663=8'd19;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd6;img686=8'd127;img687=8'd127;img688=8'd127;img689=8'd127;img690=8'd42;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd127;img715=8'd127;img716=8'd80;img717=8'd6;img718=8'd2;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd57;img148=8'd107;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd6;img158=8'd26;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd117;img176=8'd126;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd26;img186=8'd126;img187=8'd41;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd128;img204=8'd127;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd26;img214=8'd127;img215=8'd82;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd127;img232=8'd126;img233=8'd21;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd26;img242=8'd126;img243=8'd112;img244=8'd10;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd128;img260=8'd127;img261=8'd51;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd26;img270=8'd127;img271=8'd127;img272=8'd25;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd127;img288=8'd126;img289=8'd51;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd26;img298=8'd126;img299=8'd127;img300=8'd25;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd127;img316=8'd127;img317=8'd51;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd26;img326=8'd127;img327=8'd127;img328=8'd25;img329=8'd26;img330=8'd66;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd127;img344=8'd126;img345=8'd31;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd46;img354=8'd126;img355=8'd107;img356=8'd26;img357=8'd97;img358=8'd76;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd127;img372=8'd127;img373=8'd51;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd76;img382=8'd127;img383=8'd127;img384=8'd127;img385=8'd102;img386=8'd10;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd127;img400=8'd126;img401=8'd51;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd21;img409=8'd97;img410=8'd126;img411=8'd127;img412=8'd106;img413=8'd10;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd97;img428=8'd127;img429=8'd127;img430=8'd66;img431=8'd26;img432=8'd26;img433=8'd26;img434=8'd66;img435=8'd107;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd25;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd26;img456=8'd116;img457=8'd127;img458=8'd126;img459=8'd127;img460=8'd126;img461=8'd127;img462=8'd126;img463=8'd127;img464=8'd126;img465=8'd127;img466=8'd126;img467=8'd107;img468=8'd5;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd41;img485=8'd117;img486=8'd127;img487=8'd127;img488=8'd127;img489=8'd122;img490=8'd102;img491=8'd71;img492=8'd51;img493=8'd127;img494=8'd127;img495=8'd92;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd15;img514=8'd25;img515=8'd25;img516=8'd25;img517=8'd20;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd127;img522=8'd126;img523=8'd51;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd76;img550=8'd127;img551=8'd102;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd117;img578=8'd126;img579=8'd61;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd128;img606=8'd127;img607=8'd52;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd127;img634=8'd126;img635=8'd51;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd87;img662=8'd127;img663=8'd52;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd5;img690=8'd86;img691=8'd31;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd18;img101=8'd78;img102=8'd123;img103=8'd29;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd14;img128=8'd109;img129=8'd127;img130=8'd125;img131=8'd27;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd64;img156=8'd127;img157=8'd127;img158=8'd77;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd27;img183=8'd123;img184=8'd127;img185=8'd98;img186=8'd5;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd68;img211=8'd127;img212=8'd100;img213=8'd9;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd50;img238=8'd127;img239=8'd121;img240=8'd15;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd4;img265=8'd92;img266=8'd127;img267=8'd53;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd40;img293=8'd127;img294=8'd93;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd96;img320=8'd67;img321=8'd108;img322=8'd17;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd23;img347=8'd122;img348=8'd127;img349=8'd40;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd109;img375=8'd127;img376=8'd92;img377=8'd4;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd21;img382=8'd14;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd127;img403=8'd127;img404=8'd39;img405=8'd0;img406=8'd8;img407=8'd70;img408=8'd107;img409=8'd121;img410=8'd109;img411=8'd36;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd31;img430=8'd127;img431=8'd124;img432=8'd27;img433=8'd0;img434=8'd68;img435=8'd76;img436=8'd83;img437=8'd127;img438=8'd127;img439=8'd112;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd98;img458=8'd127;img459=8'd90;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd6;img465=8'd112;img466=8'd127;img467=8'd127;img468=8'd38;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd98;img486=8'd127;img487=8'd50;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd10;img493=8'd127;img494=8'd127;img495=8'd108;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd98;img514=8'd128;img515=8'd68;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd10;img521=8'd127;img522=8'd127;img523=8'd67;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd98;img542=8'd127;img543=8'd95;img544=8'd44;img545=8'd1;img546=8'd0;img547=8'd3;img548=8'd38;img549=8'd127;img550=8'd125;img551=8'd27;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd64;img570=8'd112;img571=8'd127;img572=8'd127;img573=8'd83;img574=8'd40;img575=8'd78;img576=8'd127;img577=8'd127;img578=8'd73;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd4;img598=8'd36;img599=8'd101;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd113;img606=8'd12;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd3;img628=8'd29;img629=8'd100;img630=8'd108;img631=8'd97;img632=8'd37;img633=8'd9;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd13;img173=8'd30;img174=8'd30;img175=8'd66;img176=8'd105;img177=8'd105;img178=8'd105;img179=8'd105;img180=8'd105;img181=8'd105;img182=8'd106;img183=8'd87;img184=8'd30;img185=8'd16;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd101;img201=8'd127;img202=8'd127;img203=8'd127;img204=8'd127;img205=8'd127;img206=8'd127;img207=8'd127;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd106;img214=8'd14;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd127;img229=8'd127;img230=8'd127;img231=8'd127;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd89;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd46;img257=8'd89;img258=8'd89;img259=8'd89;img260=8'd89;img261=8'd89;img262=8'd50;img263=8'd15;img264=8'd15;img265=8'd15;img266=8'd46;img267=8'd120;img268=8'd127;img269=8'd127;img270=8'd89;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd47;img295=8'd120;img296=8'd127;img297=8'd127;img298=8'd80;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd12;img321=8'd67;img322=8'd127;img323=8'd127;img324=8'd127;img325=8'd127;img326=8'd15;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd14;img345=8'd45;img346=8'd45;img347=8'd116;img348=8'd121;img349=8'd127;img350=8'd127;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd55;img355=8'd40;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd47;img372=8'd106;img373=8'd127;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd127;img383=8'd123;img384=8'd58;img385=8'd23;img386=8'd6;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd60;img400=8'd127;img401=8'd127;img402=8'd127;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd127;img413=8'd127;img414=8'd74;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd61;img428=8'd127;img429=8'd127;img430=8'd127;img431=8'd78;img432=8'd62;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd36;img438=8'd75;img439=8'd112;img440=8'd127;img441=8'd128;img442=8'd127;img443=8'd53;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd11;img456=8'd22;img457=8'd22;img458=8'd22;img459=8'd2;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd25;img468=8'd113;img469=8'd127;img470=8'd127;img471=8'd70;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd24;img497=8'd122;img498=8'd127;img499=8'd127;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd36;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd32;img525=8'd123;img526=8'd127;img527=8'd91;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd34;img541=8'd121;img542=8'd73;img543=8'd2;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd36;img552=8'd120;img553=8'd127;img554=8'd127;img555=8'd52;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd38;img569=8'd127;img570=8'd127;img571=8'd92;img572=8'd90;img573=8'd90;img574=8'd60;img575=8'd33;img576=8'd90;img577=8'd90;img578=8'd90;img579=8'd116;img580=8'd127;img581=8'd121;img582=8'd98;img583=8'd16;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd18;img597=8'd107;img598=8'd127;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd127;img607=8'd127;img608=8'd127;img609=8'd82;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd5;img626=8'd47;img627=8'd82;img628=8'd90;img629=8'd100;img630=8'd128;img631=8'd127;img632=8'd127;img633=8'd127;img634=8'd113;img635=8'd82;img636=8'd82;img637=8'd9;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd6;img657=8'd12;img658=8'd30;img659=8'd48;img660=8'd56;img661=8'd30;img662=8'd21;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd5;img164=8'd39;img165=8'd25;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd1;img187=8'd32;img188=8'd60;img189=8'd86;img190=8'd121;img191=8'd122;img192=8'd101;img193=8'd49;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd25;img210=8'd11;img211=8'd0;img212=8'd12;img213=8'd60;img214=8'd102;img215=8'd127;img216=8'd128;img217=8'd114;img218=8'd64;img219=8'd54;img220=8'd4;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd15;img236=8'd94;img237=8'd127;img238=8'd116;img239=8'd108;img240=8'd117;img241=8'd127;img242=8'd121;img243=8'd80;img244=8'd37;img245=8'd9;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd9;img263=8'd109;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd126;img268=8'd111;img269=8'd53;img270=8'd17;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd9;img290=8'd100;img291=8'd127;img292=8'd127;img293=8'd125;img294=8'd81;img295=8'd33;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd94;img318=8'd127;img319=8'd127;img320=8'd98;img321=8'd16;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd29;img345=8'd120;img346=8'd127;img347=8'd82;img348=8'd1;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd111;img373=8'd127;img374=8'd81;img375=8'd3;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd17;img400=8'd121;img401=8'd124;img402=8'd38;img403=8'd17;img404=8'd54;img405=8'd67;img406=8'd109;img407=8'd89;img408=8'd47;img409=8'd13;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd59;img428=8'd127;img429=8'd124;img430=8'd121;img431=8'd122;img432=8'd127;img433=8'd118;img434=8'd112;img435=8'd120;img436=8'd127;img437=8'd118;img438=8'd51;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd99;img456=8'd127;img457=8'd127;img458=8'd101;img459=8'd72;img460=8'd29;img461=8'd11;img462=8'd0;img463=8'd16;img464=8'd71;img465=8'd125;img466=8'd117;img467=8'd52;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd9;img484=8'd76;img485=8'd43;img486=8'd8;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd66;img494=8'd127;img495=8'd88;img496=8'd1;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd54;img522=8'd127;img523=8'd127;img524=8'd5;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd17;img549=8'd105;img550=8'd127;img551=8'd88;img552=8'd1;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd32;img576=8'd114;img577=8'd127;img578=8'd117;img579=8'd23;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd7;img601=8'd49;img602=8'd91;img603=8'd125;img604=8'd127;img605=8'd116;img606=8'd40;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd14;img623=8'd14;img624=8'd14;img625=8'd52;img626=8'd59;img627=8'd76;img628=8'd111;img629=8'd127;img630=8'd127;img631=8'd120;img632=8'd71;img633=8'd14;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd121;img651=8'd125;img652=8'd125;img653=8'd127;img654=8'd124;img655=8'd123;img656=8'd121;img657=8'd92;img658=8'd50;img659=8'd15;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd23;img680=8'd25;img681=8'd33;img682=8'd17;img683=8'd10;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd19;img127=8'd77;img128=8'd108;img129=8'd121;img130=8'd39;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd41;img154=8'd117;img155=8'd89;img156=8'd35;img157=8'd12;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd26;img177=8'd73;img178=8'd73;img179=8'd75;img180=8'd89;img181=8'd112;img182=8'd58;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd111;img205=8'd104;img206=8'd81;img207=8'd92;img208=8'd53;img209=8'd22;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd6;img232=8'd124;img233=8'd31;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd27;img260=8'd126;img261=8'd31;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd34;img288=8'd127;img289=8'd31;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd73;img316=8'd127;img317=8'd31;img318=8'd0;img319=8'd0;img320=8'd2;img321=8'd16;img322=8'd7;img323=8'd16;img324=8'd28;img325=8'd16;img326=8'd1;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd54;img344=8'd127;img345=8'd31;img346=8'd7;img347=8'd42;img348=8'd107;img349=8'd127;img350=8'd113;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd91;img355=8'd33;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd35;img372=8'd127;img373=8'd77;img374=8'd113;img375=8'd126;img376=8'd84;img377=8'd42;img378=8'd35;img379=8'd12;img380=8'd12;img381=8'd46;img382=8'd90;img383=8'd125;img384=8'd53;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd11;img400=8'd102;img401=8'd110;img402=8'd77;img403=8'd17;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd55;img412=8'd128;img413=8'd27;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd5;img440=8'd105;img441=8'd115;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd48;img469=8'd125;img470=8'd20;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd31;img497=8'd127;img498=8'd35;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd37;img525=8'd124;img526=8'd9;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd91;img553=8'd123;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd1;img569=8'd16;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd1;img579=8'd9;img580=8'd115;img581=8'd96;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd7;img597=8'd118;img598=8'd39;img599=8'd1;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd9;img606=8'd81;img607=8'd117;img608=8'd93;img609=8'd5;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd57;img626=8'd127;img627=8'd45;img628=8'd16;img629=8'd6;img630=8'd28;img631=8'd43;img632=8'd84;img633=8'd117;img634=8'd117;img635=8'd65;img636=8'd4;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd2;img654=8'd65;img655=8'd113;img656=8'd122;img657=8'd118;img658=8'd127;img659=8'd124;img660=8'd88;img661=8'd55;img662=8'd20;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd8;img94=8'd103;img95=8'd109;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd9;img121=8'd103;img122=8'd127;img123=8'd108;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd9;img148=8'd103;img149=8'd127;img150=8'd126;img151=8'd70;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd68;img176=8'd127;img177=8'd127;img178=8'd75;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd10;img203=8'd104;img204=8'd127;img205=8'd119;img206=8'd20;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd105;img231=8'd127;img232=8'd127;img233=8'd75;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd127;img259=8'd127;img260=8'd121;img261=8'd18;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd128;img287=8'd127;img288=8'd118;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd19;img297=8'd25;img298=8'd25;img299=8'd25;img300=8'd25;img301=8'd25;img302=8'd3;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd127;img315=8'd127;img316=8'd118;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd34;img323=8'd90;img324=8'd118;img325=8'd127;img326=8'd127;img327=8'd127;img328=8'd127;img329=8'd127;img330=8'd94;img331=8'd63;img332=8'd15;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd127;img343=8'd127;img344=8'd118;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd7;img350=8'd99;img351=8'd127;img352=8'd127;img353=8'd102;img354=8'd96;img355=8'd74;img356=8'd64;img357=8'd88;img358=8'd124;img359=8'd127;img360=8'd111;img361=8'd63;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd127;img371=8'd127;img372=8'd70;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd72;img378=8'd127;img379=8'd127;img380=8'd84;img381=8'd7;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd54;img387=8'd108;img388=8'd127;img389=8'd127;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd127;img399=8'd127;img400=8'd104;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd87;img406=8'd127;img407=8'd127;img408=8'd31;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd56;img416=8'd127;img417=8'd127;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd127;img427=8'd127;img428=8'd118;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd87;img434=8'd127;img435=8'd127;img436=8'd31;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd56;img444=8'd127;img445=8'd107;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd127;img455=8'd127;img456=8'd121;img457=8'd18;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd87;img462=8'd127;img463=8'd127;img464=8'd82;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd56;img472=8'd127;img473=8'd44;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd52;img483=8'd127;img484=8'd127;img485=8'd116;img486=8'd43;img487=8'd0;img488=8'd0;img489=8'd13;img490=8'd63;img491=8'd115;img492=8'd122;img493=8'd91;img494=8'd32;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd79;img500=8'd127;img501=8'd56;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd2;img511=8'd104;img512=8'd127;img513=8'd127;img514=8'd104;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd57;img520=8'd115;img521=8'd127;img522=8'd122;img523=8'd44;img524=8'd0;img525=8'd0;img526=8'd21;img527=8'd122;img528=8'd127;img529=8'd41;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd13;img540=8'd127;img541=8'd127;img542=8'd125;img543=8'd75;img544=8'd18;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd26;img549=8'd74;img550=8'd91;img551=8'd123;img552=8'd92;img553=8'd53;img554=8'd114;img555=8'd127;img556=8'd48;img557=8'd1;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd1;img568=8'd44;img569=8'd104;img570=8'd127;img571=8'd127;img572=8'd121;img573=8'd106;img574=8'd56;img575=8'd56;img576=8'd56;img577=8'd56;img578=8'd59;img579=8'd86;img580=8'd127;img581=8'd127;img582=8'd104;img583=8'd13;img584=8'd1;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd40;img598=8'd68;img599=8'd105;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd127;img607=8'd107;img608=8'd68;img609=8'd44;img610=8'd4;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd2;img628=8'd14;img629=8'd65;img630=8'd65;img631=8'd65;img632=8'd65;img633=8'd65;img634=8'd65;img635=8'd13;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd5;img152=8'd15;img153=8'd2;img154=8'd52;img155=8'd115;img156=8'd127;img157=8'd65;img158=8'd5;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd43;img180=8'd126;img181=8'd90;img182=8'd126;img183=8'd126;img184=8'd126;img185=8'd127;img186=8'd61;img187=8'd7;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd62;img208=8'd126;img209=8'd127;img210=8'd126;img211=8'd74;img212=8'd28;img213=8'd127;img214=8'd126;img215=8'd72;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd26;img235=8'd123;img236=8'd126;img237=8'd127;img238=8'd51;img239=8'd3;img240=8'd0;img241=8'd77;img242=8'd126;img243=8'd84;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd85;img263=8'd127;img264=8'd127;img265=8'd128;img266=8'd42;img267=8'd0;img268=8'd0;img269=8'd7;img270=8'd104;img271=8'd127;img272=8'd46;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd85;img291=8'd126;img292=8'd126;img293=8'd124;img294=8'd33;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd85;img299=8'd126;img300=8'd108;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd85;img319=8'd126;img320=8'd126;img321=8'd50;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd41;img327=8'd126;img328=8'd126;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd13;img346=8'd122;img347=8'd126;img348=8'd126;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd29;img355=8'd126;img356=8'd126;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd21;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd29;img383=8'd127;img384=8'd127;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd71;img402=8'd126;img403=8'd126;img404=8'd126;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd29;img411=8'd126;img412=8'd126;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd115;img430=8'd126;img431=8'd112;img432=8'd84;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd29;img439=8'd126;img440=8'd126;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd127;img458=8'd126;img459=8'd84;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd29;img467=8'd126;img468=8'd126;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd127;img486=8'd127;img487=8'd84;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd60;img495=8'd127;img496=8'd95;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd127;img514=8'd126;img515=8'd47;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd85;img523=8'd126;img524=8'd33;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd127;img542=8'd126;img543=8'd28;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd5;img550=8'd99;img551=8'd126;img552=8'd14;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd127;img570=8'd126;img571=8'd78;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd90;img578=8'd126;img579=8'd89;img580=8'd2;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd90;img598=8'd127;img599=8'd89;img600=8'd8;img601=8'd0;img602=8'd10;img603=8'd33;img604=8'd96;img605=8'd127;img606=8'd105;img607=8'd13;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd11;img626=8'd117;img627=8'd126;img628=8'd108;img629=8'd85;img630=8'd113;img631=8'd126;img632=8'd126;img633=8'd105;img634=8'd14;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd66;img655=8'd126;img656=8'd126;img657=8'd127;img658=8'd126;img659=8'd126;img660=8'd107;img661=8'd13;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd4;img683=8'd33;img684=8'd120;img685=8'd127;img686=8'd89;img687=8'd52;img688=8'd8;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd46;img149=8'd127;img150=8'd71;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd10;img176=8'd98;img177=8'd126;img178=8'd121;img179=8'd12;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd74;img189=8'd113;img190=8'd49;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd29;img204=8'd126;img205=8'd126;img206=8'd127;img207=8'd14;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd16;img216=8'd127;img217=8'd126;img218=8'd98;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd29;img232=8'd126;img233=8'd126;img234=8'd89;img235=8'd5;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd70;img244=8'd127;img245=8'd126;img246=8'd51;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd29;img260=8'd126;img261=8'd126;img262=8'd70;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd8;img271=8'd102;img272=8'd127;img273=8'd126;img274=8'd28;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd60;img288=8'd127;img289=8'd127;img290=8'd71;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd15;img299=8'd127;img300=8'd128;img301=8'd108;img302=8'd16;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd99;img316=8'd126;img317=8'd126;img318=8'd70;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd15;img327=8'd126;img328=8'd127;img329=8'd21;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd99;img344=8'd126;img345=8'd126;img346=8'd16;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd7;img354=8'd40;img355=8'd126;img356=8'd127;img357=8'd14;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd29;img371=8'd117;img372=8'd126;img373=8'd118;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd29;img382=8'd126;img383=8'd126;img384=8'd89;img385=8'd5;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd43;img399=8'd126;img400=8'd126;img401=8'd95;img402=8'd71;img403=8'd70;img404=8'd70;img405=8'd70;img406=8'd70;img407=8'd40;img408=8'd24;img409=8'd83;img410=8'd126;img411=8'd126;img412=8'd70;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd43;img427=8'd127;img428=8'd127;img429=8'd127;img430=8'd128;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd128;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd71;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd29;img455=8'd117;img456=8'd126;img457=8'd126;img458=8'd127;img459=8'd126;img460=8'd126;img461=8'd121;img462=8'd107;img463=8'd108;img464=8'd122;img465=8'd126;img466=8'd126;img467=8'd126;img468=8'd70;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd38;img484=8'd98;img485=8'd98;img486=8'd28;img487=8'd28;img488=8'd28;img489=8'd25;img490=8'd16;img491=8'd16;img492=8'd25;img493=8'd105;img494=8'd126;img495=8'd110;img496=8'd16;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd37;img521=8'd117;img522=8'd126;img523=8'd56;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd113;img549=8'd126;img550=8'd126;img551=8'd56;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd113;img577=8'd127;img578=8'd127;img579=8'd56;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd51;img604=8'd125;img605=8'd126;img606=8'd121;img607=8'd37;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd57;img632=8'd126;img633=8'd126;img634=8'd123;img635=8'd44;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd19;img660=8'd117;img661=8'd126;img662=8'd77;img663=8'd50;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd73;img689=8'd126;img690=8'd42;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd39;img156=8'd127;img157=8'd52;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd102;img184=8'd127;img185=8'd109;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd127;img212=8'd127;img213=8'd100;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd127;img240=8'd127;img241=8'd48;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd127;img268=8'd124;img269=8'd37;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd18;img295=8'd127;img296=8'd115;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd81;img323=8'd127;img324=8'd65;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd121;img351=8'd127;img352=8'd55;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd50;img378=8'd126;img379=8'd122;img380=8'd5;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd55;img406=8'd127;img407=8'd64;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd58;img434=8'd127;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd5;img461=8'd116;img462=8'd127;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd49;img489=8'd127;img490=8'd118;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd89;img517=8'd127;img518=8'd55;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd109;img545=8'd127;img546=8'd6;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd109;img573=8'd85;img574=8'd2;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd15;img600=8'd115;img601=8'd72;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd43;img628=8'd127;img629=8'd72;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd4;img656=8'd111;img657=8'd72;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd80;img685=8'd98;img686=8'd3;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd14;img210=8'd37;img211=8'd79;img212=8'd82;img213=8'd98;img214=8'd82;img215=8'd14;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd30;img236=8'd92;img237=8'd121;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd127;img243=8'd79;img244=8'd2;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd25;img262=8'd90;img263=8'd124;img264=8'd127;img265=8'd127;img266=8'd109;img267=8'd99;img268=8'd64;img269=8'd83;img270=8'd121;img271=8'd127;img272=8'd32;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd1;img288=8'd58;img289=8'd117;img290=8'd127;img291=8'd125;img292=8'd82;img293=8'd40;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd91;img299=8'd127;img300=8'd54;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd58;img316=8'd127;img317=8'd127;img318=8'd107;img319=8'd31;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd91;img327=8'd127;img328=8'd80;img329=8'd7;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd48;img343=8'd127;img344=8'd127;img345=8'd91;img346=8'd4;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd19;img354=8'd114;img355=8'd128;img356=8'd127;img357=8'd64;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd64;img371=8'd127;img372=8'd101;img373=8'd4;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd16;img380=8'd28;img381=8'd86;img382=8'd127;img383=8'd127;img384=8'd127;img385=8'd21;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd64;img399=8'd127;img400=8'd104;img401=8'd35;img402=8'd19;img403=8'd16;img404=8'd8;img405=8'd51;img406=8'd93;img407=8'd119;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd80;img413=8'd3;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd43;img427=8'd125;img428=8'd127;img429=8'd127;img430=8'd127;img431=8'd123;img432=8'd111;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd51;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd48;img456=8'd114;img457=8'd127;img458=8'd127;img459=8'd127;img460=8'd127;img461=8'd110;img462=8'd68;img463=8'd36;img464=8'd53;img465=8'd107;img466=8'd127;img467=8'd114;img468=8'd6;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd30;img486=8'd46;img487=8'd23;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd32;img493=8'd127;img494=8'd127;img495=8'd46;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd90;img521=8'd127;img522=8'd101;img523=8'd4;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd14;img548=8'd118;img549=8'd127;img550=8'd43;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd64;img576=8'd127;img577=8'd119;img578=8'd8;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd73;img604=8'd127;img605=8'd101;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd24;img631=8'd121;img632=8'd127;img633=8'd72;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd91;img659=8'd127;img660=8'd123;img661=8'd41;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd23;img686=8'd127;img687=8'd127;img688=8'd69;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd78;img714=8'd127;img715=8'd112;img716=8'd36;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd30;img742=8'd98;img743=8'd35;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd4;img191=8'd62;img192=8'd81;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd42;img217=8'd52;img218=8'd101;img219=8'd113;img220=8'd43;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd9;img241=8'd20;img242=8'd86;img243=8'd112;img244=8'd120;img245=8'd118;img246=8'd37;img247=8'd29;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd25;img266=8'd32;img267=8'd67;img268=8'd120;img269=8'd128;img270=8'd127;img271=8'd81;img272=8'd29;img273=8'd7;img274=8'd18;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd49;img291=8'd106;img292=8'd107;img293=8'd122;img294=8'd127;img295=8'd127;img296=8'd127;img297=8'd96;img298=8'd34;img299=8'd11;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd80;img319=8'd115;img320=8'd116;img321=8'd115;img322=8'd80;img323=8'd40;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd18;img346=8'd42;img347=8'd61;img348=8'd14;img349=8'd14;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd22;img373=8'd63;img374=8'd47;img375=8'd29;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd43;img401=8'd101;img402=8'd24;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd7;img429=8'd119;img430=8'd122;img431=8'd18;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd18;img457=8'd90;img458=8'd128;img459=8'd105;img460=8'd97;img461=8'd19;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd16;img486=8'd32;img487=8'd32;img488=8'd92;img489=8'd71;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd75;img517=8'd102;img518=8'd5;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd127;img545=8'd113;img546=8'd7;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd127;img573=8'd47;img574=8'd2;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd110;img601=8'd6;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd11;img627=8'd87;img628=8'd127;img629=8'd32;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd1;img654=8'd63;img655=8'd127;img656=8'd112;img657=8'd16;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd11;img682=8'd127;img683=8'd100;img684=8'd18;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd2;img710=8'd65;img711=8'd4;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd32;img199=8'd96;img200=8'd128;img201=8'd64;img202=8'd64;img203=8'd64;img204=8'd32;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd64;img227=8'd128;img228=8'd128;img229=8'd128;img230=8'd128;img231=8'd128;img232=8'd128;img233=8'd128;img234=8'd128;img235=8'd128;img236=8'd128;img237=8'd64;img238=8'd64;img239=8'd32;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd32;img255=8'd128;img256=8'd128;img257=8'd128;img258=8'd128;img259=8'd128;img260=8'd128;img261=8'd128;img262=8'd128;img263=8'd128;img264=8'd128;img265=8'd128;img266=8'd128;img267=8'd128;img268=8'd96;img269=8'd32;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd32;img285=8'd32;img286=8'd64;img287=8'd64;img288=8'd64;img289=8'd64;img290=8'd128;img291=8'd128;img292=8'd128;img293=8'd128;img294=8'd128;img295=8'd128;img296=8'd128;img297=8'd128;img298=8'd64;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd32;img322=8'd96;img323=8'd128;img324=8'd128;img325=8'd128;img326=8'd128;img327=8'd128;img328=8'd32;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd32;img352=8'd128;img353=8'd128;img354=8'd128;img355=8'd128;img356=8'd64;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd32;img381=8'd128;img382=8'd128;img383=8'd128;img384=8'd64;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd64;img410=8'd128;img411=8'd128;img412=8'd128;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd64;img438=8'd128;img439=8'd128;img440=8'd128;img441=8'd32;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd64;img466=8'd128;img467=8'd128;img468=8'd128;img469=8'd64;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd64;img494=8'd128;img495=8'd128;img496=8'd128;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd64;img522=8'd128;img523=8'd128;img524=8'd96;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd96;img550=8'd128;img551=8'd128;img552=8'd64;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd64;img577=8'd128;img578=8'd128;img579=8'd128;img580=8'd32;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd128;img605=8'd128;img606=8'd128;img607=8'd96;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd128;img633=8'd128;img634=8'd128;img635=8'd32;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd96;img660=8'd128;img661=8'd128;img662=8'd128;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd64;img687=8'd128;img688=8'd128;img689=8'd128;img690=8'd96;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd64;img715=8'd128;img716=8'd128;img717=8'd96;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd64;img743=8'd128;img744=8'd128;img745=8'd32;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd22;img154=8'd24;img155=8'd24;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd5;img180=8'd54;img181=8'd125;img182=8'd127;img183=8'd127;img184=8'd104;img185=8'd104;img186=8'd104;img187=8'd104;img188=8'd75;img189=8'd33;img190=8'd7;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd5;img207=8'd92;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd127;img216=8'd127;img217=8'd127;img218=8'd107;img219=8'd13;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd28;img234=8'd102;img235=8'd127;img236=8'd127;img237=8'd100;img238=8'd64;img239=8'd64;img240=8'd30;img241=8'd47;img242=8'd42;img243=8'd34;img244=8'd76;img245=8'd111;img246=8'd127;img247=8'd81;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd69;img262=8'd127;img263=8'd127;img264=8'd100;img265=8'd10;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd78;img274=8'd127;img275=8'd106;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd69;img290=8'd127;img291=8'd127;img292=8'd9;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd37;img301=8'd121;img302=8'd127;img303=8'd106;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd53;img318=8'd127;img319=8'd127;img320=8'd51;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd17;img328=8'd115;img329=8'd127;img330=8'd127;img331=8'd80;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd75;img347=8'd127;img348=8'd115;img349=8'd20;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd19;img354=8'd77;img355=8'd127;img356=8'd127;img357=8'd127;img358=8'd90;img359=8'd13;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd10;img375=8'd99;img376=8'd127;img377=8'd104;img378=8'd5;img379=8'd17;img380=8'd36;img381=8'd118;img382=8'd127;img383=8'd127;img384=8'd112;img385=8'd70;img386=8'd7;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd9;img404=8'd106;img405=8'd127;img406=8'd108;img407=8'd120;img408=8'd127;img409=8'd127;img410=8'd117;img411=8'd64;img412=8'd9;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd51;img432=8'd115;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd114;img437=8'd39;img438=8'd7;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd35;img457=8'd85;img458=8'd127;img459=8'd127;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd60;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd13;img482=8'd65;img483=8'd115;img484=8'd127;img485=8'd127;img486=8'd127;img487=8'd93;img488=8'd58;img489=8'd32;img490=8'd106;img491=8'd127;img492=8'd124;img493=8'd11;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd83;img509=8'd116;img510=8'd127;img511=8'd127;img512=8'd124;img513=8'd81;img514=8'd23;img515=8'd7;img516=8'd4;img517=8'd46;img518=8'd123;img519=8'd127;img520=8'd127;img521=8'd28;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd64;img537=8'd127;img538=8'd127;img539=8'd127;img540=8'd105;img541=8'd47;img542=8'd64;img543=8'd80;img544=8'd102;img545=8'd127;img546=8'd127;img547=8'd127;img548=8'd114;img549=8'd8;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd67;img566=8'd121;img567=8'd127;img568=8'd128;img569=8'd127;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd114;img576=8'd17;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd14;img595=8'd58;img596=8'd70;img597=8'd103;img598=8'd103;img599=8'd103;img600=8'd104;img601=8'd103;img602=8'd62;img603=8'd8;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd71;img179=8'd127;img180=8'd102;img181=8'd86;img182=8'd100;img183=8'd70;img184=8'd46;img185=8'd14;img186=8'd1;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd34;img206=8'd111;img207=8'd41;img208=8'd37;img209=8'd77;img210=8'd93;img211=8'd119;img212=8'd119;img213=8'd125;img214=8'd97;img215=8'd15;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd83;img234=8'd98;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd58;img242=8'd41;img243=8'd6;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd107;img262=8'd80;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd4;img289=8'd110;img290=8'd58;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd17;img317=8'd123;img318=8'd65;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd84;img346=8'd123;img347=8'd11;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd69;img353=8'd35;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd66;img374=8'd127;img375=8'd50;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd95;img381=8'd70;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd41;img402=8'd127;img403=8'd54;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd43;img408=8'd115;img409=8'd45;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd1;img430=8'd98;img431=8'd114;img432=8'd6;img433=8'd0;img434=8'd0;img435=8'd77;img436=8'd127;img437=8'd29;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd55;img459=8'd127;img460=8'd65;img461=8'd1;img462=8'd5;img463=8'd104;img464=8'd128;img465=8'd29;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd97;img488=8'd127;img489=8'd92;img490=8'd94;img491=8'd88;img492=8'd127;img493=8'd29;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd9;img516=8'd58;img517=8'd74;img518=8'd11;img519=8'd73;img520=8'd127;img521=8'd29;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd50;img548=8'd127;img549=8'd29;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd50;img576=8'd127;img577=8'd29;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd84;img604=8'd127;img605=8'd29;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd68;img632=8'd116;img633=8'd4;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd50;img660=8'd126;img661=8'd26;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd50;img688=8'd123;img689=8'd21;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd63;img716=8'd115;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd28;img96=8'd96;img97=8'd44;img98=8'd6;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd85;img124=8'd126;img125=8'd127;img126=8'd85;img127=8'd22;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd56;img152=8'd125;img153=8'd127;img154=8'd126;img155=8'd117;img156=8'd51;img157=8'd2;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd58;img181=8'd114;img182=8'd126;img183=8'd126;img184=8'd126;img185=8'd69;img186=8'd14;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd44;img210=8'd56;img211=8'd74;img212=8'd126;img213=8'd126;img214=8'd75;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd5;img240=8'd66;img241=8'd124;img242=8'd128;img243=8'd63;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd88;img270=8'd127;img271=8'd98;img272=8'd4;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd5;img298=8'd127;img299=8'd126;img300=8'd11;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd49;img326=8'd127;img327=8'd126;img328=8'd11;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd5;img352=8'd66;img353=8'd123;img354=8'd127;img355=8'd91;img356=8'd2;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd73;img374=8'd127;img375=8'd114;img376=8'd74;img377=8'd66;img378=8'd62;img379=8'd101;img380=8'd127;img381=8'd127;img382=8'd106;img383=8'd14;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd78;img402=8'd126;img403=8'd126;img404=8'd126;img405=8'd127;img406=8'd126;img407=8'd126;img408=8'd116;img409=8'd62;img410=8'd14;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd4;img430=8'd37;img431=8'd63;img432=8'd107;img433=8'd118;img434=8'd126;img435=8'd126;img436=8'd73;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd7;img462=8'd70;img463=8'd126;img464=8'd116;img465=8'd14;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd25;img491=8'd122;img492=8'd126;img493=8'd21;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd62;img512=8'd31;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd25;img519=8'd123;img520=8'd127;img521=8'd21;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd42;img539=8'd121;img540=8'd14;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd18;img545=8'd73;img546=8'd106;img547=8'd126;img548=8'd126;img549=8'd21;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd1;img566=8'd88;img567=8'd126;img568=8'd11;img569=8'd11;img570=8'd16;img571=8'd64;img572=8'd112;img573=8'd127;img574=8'd126;img575=8'd121;img576=8'd67;img577=8'd2;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd11;img594=8'd126;img595=8'd126;img596=8'd127;img597=8'd126;img598=8'd126;img599=8'd126;img600=8'd126;img601=8'd95;img602=8'd55;img603=8'd21;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd2;img622=8'd91;img623=8'd126;img624=8'd127;img625=8'd126;img626=8'd78;img627=8'd74;img628=8'd30;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd34;img201=8'd99;img202=8'd128;img203=8'd121;img204=8'd73;img205=8'd118;img206=8'd106;img207=8'd85;img208=8'd65;img209=8'd65;img210=8'd65;img211=8'd48;img212=8'd54;img213=8'd65;img214=8'd43;img215=8'd58;img216=8'd35;img217=8'd38;img218=8'd4;img219=8'd1;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd63;img229=8'd124;img230=8'd127;img231=8'd127;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd127;img243=8'd127;img244=8'd127;img245=8'd127;img246=8'd127;img247=8'd6;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd30;img258=8'd56;img259=8'd56;img260=8'd56;img261=8'd56;img262=8'd56;img263=8'd56;img264=8'd69;img265=8'd118;img266=8'd118;img267=8'd118;img268=8'd121;img269=8'd119;img270=8'd121;img271=8'd127;img272=8'd127;img273=8'd127;img274=8'd127;img275=8'd30;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd17;img297=8'd9;img298=8'd24;img299=8'd120;img300=8'd127;img301=8'd121;img302=8'd85;img303=8'd2;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd55;img327=8'd127;img328=8'd127;img329=8'd71;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd37;img354=8'd120;img355=8'd127;img356=8'd110;img357=8'd30;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd24;img374=8'd43;img375=8'd22;img376=8'd22;img377=8'd22;img378=8'd6;img379=8'd0;img380=8'd38;img381=8'd120;img382=8'd127;img383=8'd118;img384=8'd10;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd11;img401=8'd112;img402=8'd127;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd97;img407=8'd87;img408=8'd119;img409=8'd127;img410=8'd127;img411=8'd87;img412=8'd25;img413=8'd14;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd13;img429=8'd103;img430=8'd127;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd127;img441=8'd111;img442=8'd90;img443=8'd16;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd5;img458=8'd34;img459=8'd64;img460=8'd78;img461=8'd119;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd127;img466=8'd127;img467=8'd127;img468=8'd127;img469=8'd127;img470=8'd127;img471=8'd50;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd22;img489=8'd119;img490=8'd127;img491=8'd127;img492=8'd99;img493=8'd71;img494=8'd31;img495=8'd31;img496=8'd31;img497=8'd31;img498=8'd31;img499=8'd1;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd8;img516=8'd88;img517=8'd127;img518=8'd127;img519=8'd79;img520=8'd6;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd75;img544=8'd127;img545=8'd127;img546=8'd49;img547=8'd6;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd40;img571=8'd120;img572=8'd127;img573=8'd80;img574=8'd6;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd17;img598=8'd121;img599=8'd127;img600=8'd103;img601=8'd5;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd44;img626=8'd127;img627=8'd117;img628=8'd30;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd41;img653=8'd123;img654=8'd127;img655=8'd46;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd40;img680=8'd124;img681=8'd127;img682=8'd117;img683=8'd23;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd9;img707=8'd125;img708=8'd127;img709=8'd118;img710=8'd26;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd10;img735=8'd127;img736=8'd127;img737=8'd78;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd110;img157=8'd41;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd109;img185=8'd72;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd10;img208=8'd61;img209=8'd6;img210=8'd0;img211=8'd0;img212=8'd109;img213=8'd72;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd19;img236=8'd127;img237=8'd36;img238=8'd0;img239=8'd0;img240=8'd109;img241=8'd72;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd19;img264=8'd127;img265=8'd36;img266=8'd0;img267=8'd0;img268=8'd109;img269=8'd72;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd51;img292=8'd127;img293=8'd50;img294=8'd0;img295=8'd0;img296=8'd97;img297=8'd86;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd70;img320=8'd127;img321=8'd40;img322=8'd0;img323=8'd0;img324=8'd64;img325=8'd118;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd4;img347=8'd112;img348=8'd126;img349=8'd31;img350=8'd0;img351=8'd0;img352=8'd64;img353=8'd118;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd66;img375=8'd127;img376=8'd125;img377=8'd68;img378=8'd55;img379=8'd55;img380=8'd107;img381=8'd82;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd118;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd128;img407=8'd127;img408=8'd127;img409=8'd72;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd119;img431=8'd127;img432=8'd99;img433=8'd43;img434=8'd30;img435=8'd30;img436=8'd116;img437=8'd73;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd93;img459=8'd38;img460=8'd2;img461=8'd0;img462=8'd0;img463=8'd16;img464=8'd119;img465=8'd72;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd18;img492=8'd121;img493=8'd72;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd28;img520=8'd127;img521=8'd72;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd28;img548=8'd127;img549=8'd72;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd41;img576=8'd127;img577=8'd44;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd73;img604=8'd127;img605=8'd27;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd73;img632=8'd127;img633=8'd27;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd73;img660=8'd113;img661=8'd6;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd57;img688=8'd60;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd1;img68=8'd51;img69=8'd74;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd20;img96=8'd126;img97=8'd88;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd107;img124=8'd126;img125=8'd66;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd3;img150=8'd74;img151=8'd125;img152=8'd72;img153=8'd2;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd40;img178=8'd126;img179=8'd49;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd83;img206=8'd111;img207=8'd7;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd10;img216=8'd10;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd37;img233=8'd122;img234=8'd55;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd5;img242=8'd64;img243=8'd118;img244=8'd118;img245=8'd87;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd76;img261=8'd99;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd30;img269=8'd118;img270=8'd126;img271=8'd126;img272=8'd126;img273=8'd124;img274=8'd31;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd121;img289=8'd82;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd6;img296=8'd100;img297=8'd126;img298=8'd84;img299=8'd33;img300=8'd106;img301=8'd125;img302=8'd35;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd22;img316=8'd114;img317=8'd6;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd89;img324=8'd126;img325=8'd83;img326=8'd1;img327=8'd0;img328=8'd99;img329=8'd121;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd81;img344=8'd109;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd32;img351=8'd128;img352=8'd101;img353=8'd10;img354=8'd0;img355=8'd0;img356=8'd76;img357=8'd121;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd105;img372=8'd75;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd94;img379=8'd127;img380=8'd39;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd99;img385=8'd82;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd105;img400=8'd94;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd110;img407=8'd113;img408=8'd7;img409=8'd0;img410=8'd0;img411=8'd23;img412=8'd122;img413=8'd66;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd105;img428=8'd61;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd21;img434=8'd119;img435=8'd106;img436=8'd0;img437=8'd0;img438=8'd6;img439=8'd103;img440=8'd126;img441=8'd13;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd105;img456=8'd96;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd39;img462=8'd126;img463=8'd56;img464=8'd0;img465=8'd0;img466=8'd60;img467=8'd126;img468=8'd85;img469=8'd4;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd105;img484=8'd115;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd39;img490=8'd126;img491=8'd56;img492=8'd0;img493=8'd40;img494=8'd125;img495=8'd126;img496=8'd28;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd53;img512=8'd125;img513=8'd66;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd39;img518=8'd126;img519=8'd82;img520=8'd20;img521=8'd111;img522=8'd119;img523=8'd30;img524=8'd3;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd88;img541=8'd116;img542=8'd77;img543=8'd7;img544=8'd0;img545=8'd49;img546=8'd126;img547=8'd127;img548=8'd126;img549=8'd126;img550=8'd61;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd46;img569=8'd113;img570=8'd126;img571=8'd97;img572=8'd94;img573=8'd118;img574=8'd126;img575=8'd127;img576=8'd126;img577=8'd126;img578=8'd44;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd23;img598=8'd71;img599=8'd122;img600=8'd126;img601=8'd110;img602=8'd71;img603=8'd79;img604=8'd112;img605=8'd50;img606=8'd1;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd7;img161=8'd92;img162=8'd128;img163=8'd23;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd45;img188=8'd68;img189=8'd127;img190=8'd116;img191=8'd15;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd51;img215=8'd119;img216=8'd127;img217=8'd124;img218=8'd23;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd5;img233=8'd42;img234=8'd23;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd6;img242=8'd103;img243=8'd127;img244=8'd116;img245=8'd40;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd27;img260=8'd93;img261=8'd123;img262=8'd39;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd43;img270=8'd43;img271=8'd115;img272=8'd93;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd13;img287=8'd117;img288=8'd82;img289=8'd28;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd32;img298=8'd78;img299=8'd116;img300=8'd29;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd2;img313=8'd68;img314=8'd71;img315=8'd104;img316=8'd12;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd107;img326=8'd127;img327=8'd71;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd24;img341=8'd127;img342=8'd127;img343=8'd34;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd30;img353=8'd112;img354=8'd127;img355=8'd65;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd24;img369=8'd127;img370=8'd127;img371=8'd34;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd26;img381=8'd94;img382=8'd127;img383=8'd43;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd35;img397=8'd127;img398=8'd127;img399=8'd74;img400=8'd3;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd24;img408=8'd19;img409=8'd120;img410=8'd103;img411=8'd5;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd34;img425=8'd127;img426=8'd127;img427=8'd127;img428=8'd98;img429=8'd50;img430=8'd6;img431=8'd0;img432=8'd0;img433=8'd31;img434=8'd30;img435=8'd94;img436=8'd108;img437=8'd126;img438=8'd88;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd1;img453=8'd62;img454=8'd126;img455=8'd127;img456=8'd127;img457=8'd127;img458=8'd125;img459=8'd125;img460=8'd125;img461=8'd126;img462=8'd126;img463=8'd127;img464=8'd127;img465=8'd127;img466=8'd79;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd59;img483=8'd97;img484=8'd127;img485=8'd127;img486=8'd127;img487=8'd127;img488=8'd127;img489=8'd118;img490=8'd100;img491=8'd127;img492=8'd127;img493=8'd85;img494=8'd24;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd3;img512=8'd13;img513=8'd74;img514=8'd63;img515=8'd8;img516=8'd8;img517=8'd6;img518=8'd3;img519=8'd27;img520=8'd127;img521=8'd92;img522=8'd20;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd6;img548=8'd89;img549=8'd127;img550=8'd36;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd70;img576=8'd119;img577=8'd127;img578=8'd36;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd97;img604=8'd127;img605=8'd116;img606=8'd12;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd102;img632=8'd93;img633=8'd67;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd125;img660=8'd84;img661=8'd46;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd65;img688=8'd6;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd32;img149=8'd64;img150=8'd64;img151=8'd64;img152=8'd128;img153=8'd64;img154=8'd128;img155=8'd96;img156=8'd64;img157=8'd32;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd32;img176=8'd128;img177=8'd128;img178=8'd96;img179=8'd128;img180=8'd128;img181=8'd128;img182=8'd128;img183=8'd128;img184=8'd128;img185=8'd128;img186=8'd32;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd64;img204=8'd128;img205=8'd128;img206=8'd128;img207=8'd128;img208=8'd128;img209=8'd128;img210=8'd128;img211=8'd128;img212=8'd128;img213=8'd128;img214=8'd128;img215=8'd32;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd32;img232=8'd64;img233=8'd64;img234=8'd64;img235=8'd64;img236=8'd32;img237=8'd0;img238=8'd64;img239=8'd96;img240=8'd128;img241=8'd128;img242=8'd128;img243=8'd64;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd64;img268=8'd128;img269=8'd128;img270=8'd128;img271=8'd64;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd32;img293=8'd64;img294=8'd64;img295=8'd96;img296=8'd128;img297=8'd128;img298=8'd128;img299=8'd32;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd64;img320=8'd128;img321=8'd128;img322=8'd128;img323=8'd128;img324=8'd128;img325=8'd128;img326=8'd96;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd32;img347=8'd128;img348=8'd128;img349=8'd128;img350=8'd128;img351=8'd128;img352=8'd128;img353=8'd96;img354=8'd32;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd64;img374=8'd128;img375=8'd128;img376=8'd128;img377=8'd128;img378=8'd128;img379=8'd128;img380=8'd128;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd128;img402=8'd128;img403=8'd128;img404=8'd128;img405=8'd128;img406=8'd128;img407=8'd128;img408=8'd128;img409=8'd96;img410=8'd32;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd96;img430=8'd128;img431=8'd128;img432=8'd128;img433=8'd128;img434=8'd128;img435=8'd128;img436=8'd128;img437=8'd128;img438=8'd96;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd64;img459=8'd64;img460=8'd64;img461=8'd64;img462=8'd64;img463=8'd128;img464=8'd128;img465=8'd128;img466=8'd128;img467=8'd64;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd32;img492=8'd128;img493=8'd128;img494=8'd128;img495=8'd96;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd128;img521=8'd128;img522=8'd128;img523=8'd128;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd32;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd128;img549=8'd128;img550=8'd128;img551=8'd128;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd64;img571=8'd128;img572=8'd96;img573=8'd0;img574=8'd32;img575=8'd128;img576=8'd128;img577=8'd128;img578=8'd128;img579=8'd64;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd64;img598=8'd96;img599=8'd128;img600=8'd128;img601=8'd96;img602=8'd128;img603=8'd128;img604=8'd128;img605=8'd128;img606=8'd128;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd128;img627=8'd128;img628=8'd128;img629=8'd128;img630=8'd128;img631=8'd128;img632=8'd128;img633=8'd128;img634=8'd64;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd128;img655=8'd128;img656=8'd128;img657=8'd128;img658=8'd128;img659=8'd128;img660=8'd128;img661=8'd32;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd96;img684=8'd128;img685=8'd128;img686=8'd128;img687=8'd64;img688=8'd32;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd7;img153=8'd10;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd56;img180=8'd109;img181=8'd116;img182=8'd66;img183=8'd29;img184=8'd46;img185=8'd46;img186=8'd46;img187=8'd46;img188=8'd22;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd3;img206=8'd80;img207=8'd126;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd126;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd127;img216=8'd126;img217=8'd69;img218=8'd11;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd19;img233=8'd103;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd117;img240=8'd100;img241=8'd67;img242=8'd67;img243=8'd99;img244=8'd121;img245=8'd127;img246=8'd89;img247=8'd2;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd16;img260=8'd112;img261=8'd127;img262=8'd112;img263=8'd100;img264=8'd62;img265=8'd69;img266=8'd100;img267=8'd16;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd19;img273=8'd90;img274=8'd127;img275=8'd65;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd9;img287=8'd112;img288=8'd127;img289=8'd120;img290=8'd17;img291=8'd2;img292=8'd0;img293=8'd0;img294=8'd2;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd4;img302=8'd118;img303=8'd120;img304=8'd57;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd3;img314=8'd60;img315=8'd127;img316=8'd125;img317=8'd34;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd42;img331=8'd127;img332=8'd127;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd32;img342=8'd127;img343=8'd127;img344=8'd49;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd34;img359=8'd127;img360=8'd127;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd104;img370=8'd127;img371=8'd118;img372=8'd2;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd34;img387=8'd127;img388=8'd127;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd127;img398=8'd126;img399=8'd59;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd37;img415=8'd127;img416=8'd124;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd127;img426=8'd122;img427=8'd23;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd64;img443=8'd127;img444=8'd97;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd128;img454=8'd127;img455=8'd34;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd11;img470=8'd124;img471=8'd127;img472=8'd71;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd128;img482=8'd127;img483=8'd37;img484=8'd1;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd2;img496=8'd38;img497=8'd111;img498=8'd127;img499=8'd116;img500=8'd18;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd82;img510=8'd127;img511=8'd127;img512=8'd48;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd20;img522=8'd57;img523=8'd96;img524=8'd127;img525=8'd127;img526=8'd104;img527=8'd10;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd15;img538=8'd111;img539=8'd127;img540=8'd124;img541=8'd93;img542=8'd67;img543=8'd50;img544=8'd31;img545=8'd67;img546=8'd67;img547=8'd67;img548=8'd100;img549=8'd122;img550=8'd127;img551=8'd127;img552=8'd117;img553=8'd70;img554=8'd5;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd14;img567=8'd81;img568=8'd126;img569=8'd127;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd124;img579=8'd63;img580=8'd14;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd28;img597=8'd86;img598=8'd93;img599=8'd93;img600=8'd106;img601=8'd93;img602=8'd93;img603=8'd93;img604=8'd61;img605=8'd46;img606=8'd27;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd6;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd8;img207=8'd7;img208=8'd7;img209=8'd22;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd111;img227=8'd126;img228=8'd126;img229=8'd126;img230=8'd115;img231=8'd122;img232=8'd126;img233=8'd126;img234=8'd126;img235=8'd104;img236=8'd104;img237=8'd121;img238=8'd117;img239=8'd92;img240=8'd64;img241=8'd10;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd91;img255=8'd127;img256=8'd127;img257=8'd127;img258=8'd127;img259=8'd127;img260=8'd127;img261=8'd127;img262=8'd127;img263=8'd127;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd125;img270=8'd92;img271=8'd80;img272=8'd50;img273=8'd12;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd6;img284=8'd7;img285=8'd7;img286=8'd7;img287=8'd7;img288=8'd7;img289=8'd7;img290=8'd44;img291=8'd50;img292=8'd71;img293=8'd58;img294=8'd69;img295=8'd120;img296=8'd127;img297=8'd127;img298=8'd127;img299=8'd127;img300=8'd128;img301=8'd53;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd7;img324=8'd27;img325=8'd84;img326=8'd119;img327=8'd127;img328=8'd127;img329=8'd125;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd27;img355=8'd119;img356=8'd127;img357=8'd127;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd14;img383=8'd112;img384=8'd127;img385=8'd88;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd73;img411=8'd128;img412=8'd127;img413=8'd53;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd21;img438=8'd111;img439=8'd127;img440=8'd80;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd13;img465=8'd112;img466=8'd127;img467=8'd119;img468=8'd33;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd14;img492=8'd105;img493=8'd127;img494=8'd127;img495=8'd39;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd3;img519=8'd96;img520=8'd127;img521=8'd126;img522=8'd46;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd70;img547=8'd127;img548=8'd127;img549=8'd94;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd38;img574=8'd122;img575=8'd127;img576=8'd95;img577=8'd7;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd12;img601=8'd114;img602=8'd127;img603=8'd115;img604=8'd18;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd12;img628=8'd104;img629=8'd127;img630=8'd127;img631=8'd28;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd2;img655=8'd98;img656=8'd127;img657=8'd127;img658=8'd68;img659=8'd8;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd55;img683=8'd127;img684=8'd127;img685=8'd83;img686=8'd8;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd97;img711=8'd127;img712=8'd89;img713=8'd16;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd22;img739=8'd34;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd43;img124=8'd127;img125=8'd127;img126=8'd127;img127=8'd127;img128=8'd68;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd45;img151=8'd125;img152=8'd127;img153=8'd127;img154=8'd127;img155=8'd127;img156=8'd126;img157=8'd124;img158=8'd80;img159=8'd59;img160=8'd23;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd108;img179=8'd127;img180=8'd127;img181=8'd127;img182=8'd127;img183=8'd127;img184=8'd127;img185=8'd127;img186=8'd127;img187=8'd127;img188=8'd116;img189=8'd52;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd72;img206=8'd126;img207=8'd127;img208=8'd127;img209=8'd112;img210=8'd24;img211=8'd25;img212=8'd85;img213=8'd127;img214=8'd127;img215=8'd127;img216=8'd127;img217=8'd117;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd48;img233=8'd126;img234=8'd127;img235=8'd127;img236=8'd91;img237=8'd9;img238=8'd0;img239=8'd0;img240=8'd3;img241=8'd25;img242=8'd85;img243=8'd127;img244=8'd127;img245=8'd126;img246=8'd75;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd44;img260=8'd113;img261=8'd127;img262=8'd127;img263=8'd127;img264=8'd31;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd13;img271=8'd111;img272=8'd127;img273=8'd127;img274=8'd123;img275=8'd21;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd20;img287=8'd123;img288=8'd127;img289=8'd127;img290=8'd127;img291=8'd69;img292=8'd4;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd21;img300=8'd111;img301=8'd127;img302=8'd127;img303=8'd59;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd59;img315=8'd127;img316=8'd127;img317=8'd127;img318=8'd113;img319=8'd14;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd78;img329=8'd127;img330=8'd127;img331=8'd59;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd59;img343=8'd127;img344=8'd127;img345=8'd127;img346=8'd29;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd78;img357=8'd127;img358=8'd127;img359=8'd59;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd76;img371=8'd127;img372=8'd127;img373=8'd89;img374=8'd4;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd78;img385=8'd127;img386=8'd127;img387=8'd109;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd124;img399=8'd127;img400=8'd127;img401=8'd29;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd78;img413=8'd127;img414=8'd127;img415=8'd124;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd77;img427=8'd127;img428=8'd127;img429=8'd60;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd78;img441=8'd127;img442=8'd127;img443=8'd110;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd104;img455=8'd127;img456=8'd127;img457=8'd78;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd0;img467=8'd3;img468=8'd87;img469=8'd127;img470=8'd127;img471=8'd59;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd80;img483=8'd127;img484=8'd127;img485=8'd78;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd4;img495=8'd67;img496=8'd127;img497=8'd127;img498=8'd127;img499=8'd59;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd59;img511=8'd127;img512=8'd127;img513=8'd78;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd3;img522=8'd34;img523=8'd127;img524=8'd127;img525=8'd127;img526=8'd126;img527=8'd51;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd23;img539=8'd123;img540=8'd127;img541=8'd108;img542=8'd17;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd4;img548=8'd14;img549=8'd67;img550=8'd127;img551=8'd127;img552=8'd127;img553=8'd126;img554=8'd74;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd121;img568=8'd127;img569=8'd127;img570=8'd108;img571=8'd20;img572=8'd64;img573=8'd75;img574=8'd75;img575=8'd87;img576=8'd127;img577=8'd127;img578=8'd127;img579=8'd127;img580=8'd126;img581=8'd108;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd53;img596=8'd122;img597=8'd127;img598=8'd127;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd127;img607=8'd127;img608=8'd77;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd115;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd125;img629=8'd127;img630=8'd127;img631=8'd111;img632=8'd105;img633=8'd78;img634=8'd92;img635=8'd59;img636=8'd23;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd81;img654=8'd70;img655=8'd117;img656=8'd42;img657=8'd62;img658=8'd62;img659=8'd48;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd24;img120=8'd68;img121=8'd121;img122=8'd127;img123=8'd127;img124=8'd127;img125=8'd127;img126=8'd127;img127=8'd128;img128=8'd101;img129=8'd65;img130=8'd4;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd17;img147=8'd114;img148=8'd127;img149=8'd127;img150=8'd127;img151=8'd127;img152=8'd116;img153=8'd68;img154=8'd96;img155=8'd109;img156=8'd117;img157=8'd127;img158=8'd98;img159=8'd27;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd22;img175=8'd120;img176=8'd127;img177=8'd127;img178=8'd126;img179=8'd95;img180=8'd16;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd19;img185=8'd73;img186=8'd127;img187=8'd89;img188=8'd8;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd41;img204=8'd91;img205=8'd91;img206=8'd34;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd2;img214=8'd71;img215=8'd127;img216=8'd79;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd3;img243=8'd91;img244=8'd121;img245=8'd43;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd59;img272=8'd127;img273=8'd85;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd24;img300=8'd127;img301=8'd85;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd24;img328=8'd127;img329=8'd85;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd62;img356=8'd127;img357=8'd85;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd83;img384=8'd127;img385=8'd44;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd5;img411=8'd96;img412=8'd102;img413=8'd6;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd3;img438=8'd57;img439=8'd127;img440=8'd94;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd6;img466=8'd127;img467=8'd127;img468=8'd41;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd2;img484=8'd27;img485=8'd65;img486=8'd9;img487=8'd3;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd3;img493=8'd95;img494=8'd127;img495=8'd73;img496=8'd1;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd16;img511=8'd89;img512=8'd127;img513=8'd127;img514=8'd127;img515=8'd97;img516=8'd74;img517=8'd61;img518=8'd4;img519=8'd0;img520=8'd64;img521=8'd127;img522=8'd118;img523=8'd19;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd12;img538=8'd92;img539=8'd127;img540=8'd108;img541=8'd51;img542=8'd101;img543=8'd105;img544=8'd127;img545=8'd127;img546=8'd93;img547=8'd83;img548=8'd123;img549=8'd126;img550=8'd64;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd18;img566=8'd127;img567=8'd101;img568=8'd7;img569=8'd0;img570=8'd0;img571=8'd4;img572=8'd45;img573=8'd117;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd121;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd18;img594=8'd127;img595=8'd120;img596=8'd53;img597=8'd5;img598=8'd0;img599=8'd24;img600=8'd79;img601=8'd119;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd126;img606=8'd66;img607=8'd15;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd11;img622=8'd87;img623=8'd127;img624=8'd127;img625=8'd112;img626=8'd110;img627=8'd119;img628=8'd127;img629=8'd127;img630=8'd112;img631=8'd27;img632=8'd44;img633=8'd126;img634=8'd127;img635=8'd67;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd2;img651=8'd25;img652=8'd116;img653=8'd127;img654=8'd127;img655=8'd127;img656=8'd117;img657=8'd54;img658=8'd6;img659=8'd0;img660=8'd0;img661=8'd42;img662=8'd127;img663=8'd125;img664=8'd61;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd23;img181=8'd77;img182=8'd104;img183=8'd124;img184=8'd115;img185=8'd127;img186=8'd128;img187=8'd69;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd20;img208=8'd103;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd107;img216=8'd16;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd9;img235=8'd105;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd118;img241=8'd127;img242=8'd127;img243=8'd127;img244=8'd63;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd49;img263=8'd127;img264=8'd127;img265=8'd127;img266=8'd76;img267=8'd20;img268=8'd13;img269=8'd76;img270=8'd127;img271=8'd127;img272=8'd84;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd83;img291=8'd127;img292=8'd127;img293=8'd101;img294=8'd22;img295=8'd0;img296=8'd5;img297=8'd104;img298=8'd127;img299=8'd127;img300=8'd103;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd27;img319=8'd126;img320=8'd127;img321=8'd121;img322=8'd42;img323=8'd68;img324=8'd90;img325=8'd127;img326=8'd127;img327=8'd127;img328=8'd63;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd95;img348=8'd127;img349=8'd127;img350=8'd127;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd127;img355=8'd127;img356=8'd32;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd2;img376=8'd28;img377=8'd105;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd127;img383=8'd101;img384=8'd1;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd44;img406=8'd114;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd119;img411=8'd46;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd52;img434=8'd124;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd31;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd46;img461=8'd124;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd83;img466=8'd1;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd50;img488=8'd115;img489=8'd127;img490=8'd127;img491=8'd85;img492=8'd57;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd48;img515=8'd127;img516=8'd127;img517=8'd127;img518=8'd115;img519=8'd8;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd48;img542=8'd114;img543=8'd127;img544=8'd127;img545=8'd127;img546=8'd67;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd19;img569=8'd114;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd101;img574=8'd10;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd97;img597=8'd127;img598=8'd127;img599=8'd127;img600=8'd101;img601=8'd11;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd46;img624=8'd123;img625=8'd127;img626=8'd127;img627=8'd121;img628=8'd45;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd18;img651=8'd121;img652=8'd127;img653=8'd127;img654=8'd127;img655=8'd71;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd107;img680=8'd127;img681=8'd127;img682=8'd93;img683=8'd12;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd92;img708=8'd127;img709=8'd124;img710=8'd12;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd12;img153=8'd110;img154=8'd128;img155=8'd53;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd21;img181=8'd127;img182=8'd127;img183=8'd79;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd34;img209=8'd127;img210=8'd127;img211=8'd79;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd80;img237=8'd127;img238=8'd127;img239=8'd79;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd80;img265=8'd127;img266=8'd127;img267=8'd79;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd80;img293=8'd127;img294=8'd127;img295=8'd79;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd80;img321=8'd127;img322=8'd127;img323=8'd79;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd80;img349=8'd127;img350=8'd127;img351=8'd79;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd43;img377=8'd127;img378=8'd127;img379=8'd109;img380=8'd8;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd21;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd12;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd21;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd12;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd21;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd12;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd21;img489=8'd127;img490=8'd127;img491=8'd127;img492=8'd12;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd21;img517=8'd127;img518=8'd127;img519=8'd103;img520=8'd6;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd21;img545=8'd127;img546=8'd127;img547=8'd79;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd32;img573=8'd127;img574=8'd127;img575=8'd79;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd6;img600=8'd102;img601=8'd127;img602=8'd127;img603=8'd37;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd80;img629=8'd127;img630=8'd96;img631=8'd5;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd11;img656=8'd121;img657=8'd127;img658=8'd88;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd1;img684=8'd56;img685=8'd85;img686=8'd75;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd19;img214=8'd113;img215=8'd107;img216=8'd10;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd7;img229=8'd13;img230=8'd13;img231=8'd10;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd6;img236=8'd13;img237=8'd7;img238=8'd13;img239=8'd13;img240=8'd24;img241=8'd112;img242=8'd127;img243=8'd123;img244=8'd16;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd73;img257=8'd127;img258=8'd127;img259=8'd115;img260=8'd33;img261=8'd68;img262=8'd79;img263=8'd100;img264=8'd127;img265=8'd105;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd127;img270=8'd127;img271=8'd76;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd59;img285=8'd106;img286=8'd111;img287=8'd103;img288=8'd110;img289=8'd115;img290=8'd127;img291=8'd127;img292=8'd127;img293=8'd127;img294=8'd127;img295=8'd127;img296=8'd127;img297=8'd127;img298=8'd91;img299=8'd8;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd6;img314=8'd12;img315=8'd0;img316=8'd11;img317=8'd19;img318=8'd36;img319=8'd36;img320=8'd36;img321=8'd36;img322=8'd36;img323=8'd92;img324=8'd127;img325=8'd120;img326=8'd23;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd4;img351=8'd93;img352=8'd127;img353=8'd51;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd62;img379=8'd127;img380=8'd127;img381=8'd36;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd73;img407=8'd127;img408=8'd118;img409=8'd23;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd48;img431=8'd55;img432=8'd55;img433=8'd55;img434=8'd96;img435=8'd127;img436=8'd125;img437=8'd72;img438=8'd55;img439=8'd55;img440=8'd84;img441=8'd32;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd41;img458=8'd126;img459=8'd127;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd127;img466=8'd127;img467=8'd127;img468=8'd127;img469=8'd44;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd53;img487=8'd116;img488=8'd121;img489=8'd122;img490=8'd127;img491=8'd127;img492=8'd123;img493=8'd92;img494=8'd75;img495=8'd41;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd7;img518=8'd127;img519=8'd125;img520=8'd38;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd7;img546=8'd127;img547=8'd109;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd47;img574=8'd127;img575=8'd109;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd67;img602=8'd127;img603=8'd109;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd113;img630=8'd127;img631=8'd91;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd127;img658=8'd127;img659=8'd48;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd127;img686=8'd127;img687=8'd48;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd127;img714=8'd127;img715=8'd48;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd41;img742=8'd121;img743=8'd26;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd27;img125=8'd88;img126=8'd115;img127=8'd127;img128=8'd66;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd33;img152=8'd118;img153=8'd105;img154=8'd123;img155=8'd127;img156=8'd121;img157=8'd30;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd21;img179=8'd118;img180=8'd103;img181=8'd27;img182=8'd17;img183=8'd74;img184=8'd127;img185=8'd75;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd91;img207=8'd109;img208=8'd4;img209=8'd0;img210=8'd0;img211=8'd16;img212=8'd121;img213=8'd57;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd36;img235=8'd53;img236=8'd1;img237=8'd0;img238=8'd0;img239=8'd16;img240=8'd118;img241=8'd38;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd8;img267=8'd80;img268=8'd111;img269=8'd40;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd5;img294=8'd108;img295=8'd127;img296=8'd76;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd31;img321=8'd109;img322=8'd127;img323=8'd87;img324=8'd12;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd4;img347=8'd72;img348=8'd125;img349=8'd127;img350=8'd123;img351=8'd22;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd66;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd96;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd23;img403=8'd112;img404=8'd120;img405=8'd82;img406=8'd115;img407=8'd76;img408=8'd88;img409=8'd63;img410=8'd1;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd14;img436=8'd114;img437=8'd127;img438=8'd85;img439=8'd23;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd5;img465=8'd74;img466=8'd127;img467=8'd67;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd4;img494=8'd110;img495=8'd90;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd92;img523=8'd120;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd32;img550=8'd127;img551=8'd77;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd18;img569=8'd5;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd2;img576=8'd44;img577=8'd104;img578=8'd127;img579=8'd10;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd6;img596=8'd81;img597=8'd60;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd2;img603=8'd74;img604=8'd127;img605=8'd127;img606=8'd87;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd14;img624=8'd123;img625=8'd104;img626=8'd18;img627=8'd6;img628=8'd12;img629=8'd45;img630=8'd113;img631=8'd127;img632=8'd127;img633=8'd99;img634=8'd9;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd95;img653=8'd128;img654=8'd124;img655=8'd121;img656=8'd122;img657=8'd127;img658=8'd128;img659=8'd117;img660=8'd40;img661=8'd4;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd2;img206=8'd19;img207=8'd64;img208=8'd70;img209=8'd70;img210=8'd70;img211=8'd29;img212=8'd8;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd24;img232=8'd59;img233=8'd97;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd108;img241=8'd40;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd51;img259=8'd99;img260=8'd127;img261=8'd115;img262=8'd78;img263=8'd17;img264=8'd10;img265=8'd10;img266=8'd21;img267=8'd62;img268=8'd126;img269=8'd124;img270=8'd81;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd32;img286=8'd118;img287=8'd122;img288=8'd53;img289=8'd3;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd53;img297=8'd127;img298=8'd122;img299=8'd26;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd121;img314=8'd127;img315=8'd63;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd3;img325=8'd100;img326=8'd127;img327=8'd36;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd128;img342=8'd127;img343=8'd57;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd96;img354=8'd127;img355=8'd36;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd52;img370=8'd32;img371=8'd10;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd18;img381=8'd122;img382=8'd114;img383=8'd6;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd64;img409=8'd127;img410=8'd69;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd60;img436=8'd127;img437=8'd71;img438=8'd2;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd35;img463=8'd127;img464=8'd107;img465=8'd14;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd60;img490=8'd115;img491=8'd92;img492=8'd14;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd11;img516=8'd80;img517=8'd125;img518=8'd90;img519=8'd2;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd97;img544=8'd127;img545=8'd104;img546=8'd40;img547=8'd8;img548=8'd16;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd9;img556=8'd24;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd7;img570=8'd77;img571=8'd125;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd117;img576=8'd118;img577=8'd112;img578=8'd114;img579=8'd114;img580=8'd114;img581=8'd101;img582=8'd65;img583=8'd117;img584=8'd122;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd35;img598=8'd127;img599=8'd65;img600=8'd42;img601=8'd42;img602=8'd42;img603=8'd42;img604=8'd35;img605=8'd71;img606=8'd72;img607=8'd77;img608=8'd46;img609=8'd107;img610=8'd72;img611=8'd115;img612=8'd127;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd2;img626=8'd18;img627=8'd10;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd8;img638=8'd0;img639=8'd12;img640=8'd18;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd35;img184=8'd101;img185=8'd128;img186=8'd63;img187=8'd1;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd36;img211=8'd120;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd5;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd9;img238=8'd121;img239=8'd127;img240=8'd97;img241=8'd83;img242=8'd127;img243=8'd7;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd26;img265=8'd101;img266=8'd127;img267=8'd90;img268=8'd4;img269=8'd30;img270=8'd127;img271=8'd60;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd36;img292=8'd106;img293=8'd124;img294=8'd52;img295=8'd7;img296=8'd0;img297=8'd30;img298=8'd127;img299=8'd77;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd33;img319=8'd122;img320=8'd125;img321=8'd67;img322=8'd0;img323=8'd5;img324=8'd62;img325=8'd117;img326=8'd127;img327=8'd88;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd8;img346=8'd116;img347=8'd127;img348=8'd73;img349=8'd26;img350=8'd79;img351=8'd117;img352=8'd127;img353=8'd127;img354=8'd127;img355=8'd26;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd27;img374=8'd123;img375=8'd127;img376=8'd104;img377=8'd125;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd110;img383=8'd4;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd110;img403=8'd127;img404=8'd127;img405=8'd120;img406=8'd127;img407=8'd127;img408=8'd126;img409=8'd93;img410=8'd7;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd22;img431=8'd46;img432=8'd46;img433=8'd24;img434=8'd127;img435=8'd127;img436=8'd70;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd82;img462=8'd127;img463=8'd71;img464=8'd2;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd41;img489=8'd126;img490=8'd127;img491=8'd27;img492=8'd0;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd79;img517=8'd127;img518=8'd109;img519=8'd9;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd20;img544=8'd121;img545=8'd124;img546=8'd39;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd77;img572=8'd127;img573=8'd113;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd4;img599=8'd112;img600=8'd127;img601=8'd51;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd6;img627=8'd127;img628=8'd127;img629=8'd11;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd59;img655=8'd127;img656=8'd127;img657=8'd29;img658=8'd59;img659=8'd27;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd22;img683=8'd127;img684=8'd127;img685=8'd127;img686=8'd119;img687=8'd20;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd1;img711=8'd86;img712=8'd127;img713=8'd100;img714=8'd34;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd16;img210=8'd59;img211=8'd104;img212=8'd127;img213=8'd127;img214=8'd127;img215=8'd128;img216=8'd127;img217=8'd69;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd37;img232=8'd58;img233=8'd117;img234=8'd117;img235=8'd117;img236=8'd117;img237=8'd120;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd127;img243=8'd127;img244=8'd127;img245=8'd114;img246=8'd19;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd15;img258=8'd96;img259=8'd122;img260=8'd127;img261=8'd127;img262=8'd127;img263=8'd127;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd127;img270=8'd127;img271=8'd127;img272=8'd127;img273=8'd127;img274=8'd48;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd49;img286=8'd127;img287=8'd127;img288=8'd127;img289=8'd127;img290=8'd127;img291=8'd127;img292=8'd127;img293=8'd127;img294=8'd127;img295=8'd127;img296=8'd127;img297=8'd127;img298=8'd127;img299=8'd127;img300=8'd127;img301=8'd111;img302=8'd12;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd42;img314=8'd124;img315=8'd127;img316=8'd127;img317=8'd127;img318=8'd127;img319=8'd127;img320=8'd127;img321=8'd122;img322=8'd110;img323=8'd110;img324=8'd73;img325=8'd127;img326=8'd127;img327=8'd127;img328=8'd127;img329=8'd106;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd43;img343=8'd66;img344=8'd111;img345=8'd52;img346=8'd52;img347=8'd52;img348=8'd52;img349=8'd38;img350=8'd0;img351=8'd0;img352=8'd8;img353=8'd127;img354=8'd127;img355=8'd127;img356=8'd127;img357=8'd106;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd43;img380=8'd100;img381=8'd127;img382=8'd127;img383=8'd127;img384=8'd127;img385=8'd71;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd11;img407=8'd102;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd67;img413=8'd1;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd13;img434=8'd98;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd27;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd13;img461=8'd97;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd127;img466=8'd113;img467=8'd70;img468=8'd5;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd95;img489=8'd127;img490=8'd127;img491=8'd127;img492=8'd127;img493=8'd115;img494=8'd24;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd44;img516=8'd122;img517=8'd127;img518=8'd127;img519=8'd127;img520=8'd125;img521=8'd23;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd4;img542=8'd72;img543=8'd126;img544=8'd127;img545=8'd127;img546=8'd127;img547=8'd125;img548=8'd83;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd41;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd45;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd45;img597=8'd124;img598=8'd127;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd76;img603=8'd3;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd47;img624=8'd122;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd127;img629=8'd97;img630=8'd5;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd96;img652=8'd127;img653=8'd127;img654=8'd127;img655=8'd127;img656=8'd116;img657=8'd33;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd44;img680=8'd120;img681=8'd127;img682=8'd127;img683=8'd127;img684=8'd106;img685=8'd13;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd81;img709=8'd127;img710=8'd127;img711=8'd127;img712=8'd39;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd8;img737=8'd62;img738=8'd127;img739=8'd60;img740=8'd6;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd62;img206=8'd87;img207=8'd26;img208=8'd7;img209=8'd0;img210=8'd4;img211=8'd39;img212=8'd118;img213=8'd25;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd127;img234=8'd126;img235=8'd126;img236=8'd106;img237=8'd95;img238=8'd101;img239=8'd126;img240=8'd126;img241=8'd82;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd127;img262=8'd126;img263=8'd126;img264=8'd126;img265=8'd126;img266=8'd127;img267=8'd126;img268=8'd126;img269=8'd124;img270=8'd19;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd36;img289=8'd127;img290=8'd126;img291=8'd49;img292=8'd77;img293=8'd108;img294=8'd127;img295=8'd126;img296=8'd126;img297=8'd126;img298=8'd21;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd53;img317=8'd127;img318=8'd126;img319=8'd11;img320=8'd0;img321=8'd9;img322=8'd21;img323=8'd21;img324=8'd118;img325=8'd126;img326=8'd21;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd54;img345=8'd128;img346=8'd127;img347=8'd11;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd117;img353=8'd127;img354=8'd30;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd53;img373=8'd127;img374=8'd126;img375=8'd11;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd116;img381=8'd126;img382=8'd74;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd53;img401=8'd127;img402=8'd126;img403=8'd11;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd116;img409=8'd126;img410=8'd74;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd40;img429=8'd114;img430=8'd126;img431=8'd11;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd116;img437=8'd126;img438=8'd74;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd21;img458=8'd74;img459=8'd6;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd116;img465=8'd126;img466=8'd74;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd117;img493=8'd127;img494=8'd74;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd116;img521=8'd126;img522=8'd74;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd116;img549=8'd126;img550=8'd74;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd116;img577=8'd126;img578=8'd74;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd116;img605=8'd126;img606=8'd74;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd117;img633=8'd127;img634=8'd105;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd116;img661=8'd126;img662=8'd126;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd116;img689=8'd126;img690=8'd126;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd116;img717=8'd126;img718=8'd126;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd24;img745=8'd109;img746=8'd82;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd40;img100=8'd84;img101=8'd70;img102=8'd2;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd41;img126=8'd99;img127=8'd122;img128=8'd127;img129=8'd127;img130=8'd8;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd2;img152=8'd44;img153=8'd127;img154=8'd127;img155=8'd127;img156=8'd127;img157=8'd127;img158=8'd8;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd25;img180=8'd127;img181=8'd127;img182=8'd127;img183=8'd127;img184=8'd104;img185=8'd67;img186=8'd2;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd4;img207=8'd88;img208=8'd127;img209=8'd127;img210=8'd119;img211=8'd53;img212=8'd5;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd73;img235=8'd128;img236=8'd127;img237=8'd126;img238=8'd15;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd10;img262=8'd107;img263=8'd127;img264=8'd113;img265=8'd24;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd100;img290=8'd127;img291=8'd126;img292=8'd52;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd118;img318=8'd128;img319=8'd76;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd118;img346=8'd127;img347=8'd67;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd34;img373=8'd126;img374=8'd113;img375=8'd20;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd9;img381=8'd50;img382=8'd99;img383=8'd86;img384=8'd5;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd35;img401=8'd126;img402=8'd91;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd38;img408=8'd125;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd52;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd118;img430=8'd91;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd10;img435=8'd111;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd117;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd118;img458=8'd91;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd54;img463=8'd127;img464=8'd127;img465=8'd122;img466=8'd84;img467=8'd108;img468=8'd117;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd118;img486=8'd102;img487=8'd5;img488=8'd0;img489=8'd1;img490=8'd93;img491=8'd127;img492=8'd121;img493=8'd37;img494=8'd5;img495=8'd103;img496=8'd117;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd113;img514=8'd128;img515=8'd67;img516=8'd4;img517=8'd3;img518=8'd127;img519=8'd127;img520=8'd60;img521=8'd0;img522=8'd46;img523=8'd127;img524=8'd87;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd52;img542=8'd127;img543=8'd127;img544=8'd88;img545=8'd36;img546=8'd127;img547=8'd127;img548=8'd74;img549=8'd53;img550=8'd125;img551=8'd127;img552=8'd13;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd2;img570=8'd91;img571=8'd127;img572=8'd127;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd127;img579=8'd92;img580=8'd2;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd67;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd117;img606=8'd92;img607=8'd14;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd2;img628=8'd36;img629=8'd119;img630=8'd117;img631=8'd75;img632=8'd67;img633=8'd15;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd1;img97=8'd9;img98=8'd9;img99=8'd28;img100=8'd69;img101=8'd96;img102=8'd66;img103=8'd4;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd8;img123=8'd48;img124=8'd82;img125=8'd127;img126=8'd127;img127=8'd127;img128=8'd127;img129=8'd127;img130=8'd127;img131=8'd89;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd21;img149=8'd76;img150=8'd104;img151=8'd127;img152=8'd127;img153=8'd127;img154=8'd127;img155=8'd127;img156=8'd127;img157=8'd127;img158=8'd127;img159=8'd113;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd95;img177=8'd127;img178=8'd127;img179=8'd127;img180=8'd127;img181=8'd105;img182=8'd78;img183=8'd33;img184=8'd33;img185=8'd74;img186=8'd127;img187=8'd124;img188=8'd33;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd35;img205=8'd119;img206=8'd127;img207=8'd83;img208=8'd24;img209=8'd9;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd57;img214=8'd127;img215=8'd127;img216=8'd45;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd12;img234=8'd15;img235=8'd1;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd57;img242=8'd127;img243=8'd127;img244=8'd45;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd4;img270=8'd125;img271=8'd127;img272=8'd45;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd57;img298=8'd127;img299=8'd127;img300=8'd45;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd94;img326=8'd127;img327=8'd125;img328=8'd37;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd34;img353=8'd124;img354=8'd127;img355=8'd113;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd94;img381=8'd127;img382=8'd126;img383=8'd51;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd15;img408=8'd115;img409=8'd127;img410=8'd122;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd14;img435=8'd106;img436=8'd127;img437=8'd127;img438=8'd122;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd2;img456=8'd23;img457=8'd114;img458=8'd125;img459=8'd125;img460=8'd125;img461=8'd125;img462=8'd126;img463=8'd127;img464=8'd127;img465=8'd127;img466=8'd33;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd34;img484=8'd127;img485=8'd127;img486=8'd127;img487=8'd127;img488=8'd127;img489=8'd127;img490=8'd128;img491=8'd127;img492=8'd127;img493=8'd127;img494=8'd73;img495=8'd14;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd23;img511=8'd113;img512=8'd127;img513=8'd127;img514=8'd127;img515=8'd127;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd127;img520=8'd127;img521=8'd127;img522=8'd127;img523=8'd122;img524=8'd40;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd77;img539=8'd127;img540=8'd127;img541=8'd127;img542=8'd127;img543=8'd127;img544=8'd127;img545=8'd127;img546=8'd120;img547=8'd49;img548=8'd85;img549=8'd109;img550=8'd127;img551=8'd127;img552=8'd121;img553=8'd77;img554=8'd7;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd77;img567=8'd127;img568=8'd127;img569=8'd127;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd91;img574=8'd21;img575=8'd0;img576=8'd0;img577=8'd12;img578=8'd57;img579=8'd110;img580=8'd127;img581=8'd127;img582=8'd87;img583=8'd6;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd77;img595=8'd127;img596=8'd127;img597=8'd127;img598=8'd127;img599=8'd126;img600=8'd44;img601=8'd7;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd11;img608=8'd29;img609=8'd90;img610=8'd127;img611=8'd41;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd14;img623=8'd108;img624=8'd127;img625=8'd127;img626=8'd75;img627=8'd11;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd18;img638=8'd68;img639=8'd41;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd46;img205=8'd94;img206=8'd32;img207=8'd20;img208=8'd15;img209=8'd0;img210=8'd9;img211=8'd0;img212=8'd9;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd98;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd120;img237=8'd93;img238=8'd108;img239=8'd93;img240=8'd108;img241=8'd93;img242=8'd93;img243=8'd16;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd60;img261=8'd127;img262=8'd107;img263=8'd120;img264=8'd113;img265=8'd90;img266=8'd125;img267=8'd125;img268=8'd125;img269=8'd127;img270=8'd127;img271=8'd69;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd93;img289=8'd127;img290=8'd30;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd123;img298=8'd127;img299=8'd76;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd31;img316=8'd124;img317=8'd92;img318=8'd8;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd37;img325=8'd126;img326=8'd127;img327=8'd35;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd11;img343=8'd105;img344=8'd125;img345=8'd26;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd50;img353=8'd127;img354=8'd127;img355=8'd22;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd46;img371=8'd127;img372=8'd88;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd60;img381=8'd127;img382=8'd121;img383=8'd18;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd6;img399=8'd47;img400=8'd22;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd104;img409=8'd127;img410=8'd95;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd104;img437=8'd127;img438=8'd91;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd104;img465=8'd127;img466=8'd41;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd104;img493=8'd127;img494=8'd41;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd104;img521=8'd127;img522=8'd41;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd8;img548=8'd109;img549=8'd124;img550=8'd31;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd30;img576=8'd127;img577=8'd114;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd82;img604=8'd127;img605=8'd114;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd84;img632=8'd127;img633=8'd114;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd84;img660=8'd127;img661=8'd114;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd7;img687=8'd108;img688=8'd127;img689=8'd84;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd11;img715=8'd127;img716=8'd127;img717=8'd60;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd2;img743=8'd91;img744=8'd107;img745=8'd11;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd3;img157=8'd38;img158=8'd0;img159=8'd49;img160=8'd93;img161=8'd89;img162=8'd47;img163=8'd10;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd8;img182=8'd56;img183=8'd98;img184=8'd119;img185=8'd47;img186=8'd0;img187=8'd104;img188=8'd125;img189=8'd127;img190=8'd127;img191=8'd58;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd10;img207=8'd25;img208=8'd54;img209=8'd99;img210=8'd123;img211=8'd92;img212=8'd13;img213=8'd0;img214=8'd0;img215=8'd41;img216=8'd123;img217=8'd127;img218=8'd125;img219=8'd46;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd9;img233=8'd42;img234=8'd115;img235=8'd127;img236=8'd127;img237=8'd111;img238=8'd43;img239=8'd0;img240=8'd0;img241=8'd1;img242=8'd63;img243=8'd127;img244=8'd127;img245=8'd89;img246=8'd27;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd67;img261=8'd127;img262=8'd127;img263=8'd109;img264=8'd59;img265=8'd2;img266=8'd0;img267=8'd0;img268=8'd31;img269=8'd101;img270=8'd127;img271=8'd121;img272=8'd66;img273=8'd4;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd54;img288=8'd122;img289=8'd127;img290=8'd107;img291=8'd23;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd31;img296=8'd120;img297=8'd127;img298=8'd110;img299=8'd15;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd22;img315=8'd123;img316=8'd127;img317=8'd105;img318=8'd25;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd16;img323=8'd121;img324=8'd127;img325=8'd111;img326=8'd14;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd48;img343=8'd127;img344=8'd127;img345=8'd28;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd9;img350=8'd99;img351=8'd127;img352=8'd109;img353=8'd14;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd14;img371=8'd110;img372=8'd127;img373=8'd117;img374=8'd72;img375=8'd20;img376=8'd21;img377=8'd102;img378=8'd127;img379=8'd103;img380=8'd5;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd58;img400=8'd124;img401=8'd127;img402=8'd127;img403=8'd122;img404=8'd117;img405=8'd127;img406=8'd112;img407=8'd12;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd19;img429=8'd42;img430=8'd84;img431=8'd123;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd104;img436=8'd58;img437=8'd5;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd7;img459=8'd118;img460=8'd127;img461=8'd115;img462=8'd82;img463=8'd119;img464=8'd122;img465=8'd106;img466=8'd40;img467=8'd1;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd50;img487=8'd127;img488=8'd127;img489=8'd50;img490=8'd0;img491=8'd0;img492=8'd19;img493=8'd113;img494=8'd127;img495=8'd65;img496=8'd4;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd36;img515=8'd127;img516=8'd115;img517=8'd6;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd1;img522=8'd85;img523=8'd127;img524=8'd26;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd48;img543=8'd127;img544=8'd127;img545=8'd9;img546=8'd0;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd41;img551=8'd127;img552=8'd99;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd40;img571=8'd127;img572=8'd127;img573=8'd9;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd66;img579=8'd127;img580=8'd60;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd3;img599=8'd107;img600=8'd127;img601=8'd39;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd1;img606=8'd92;img607=8'd122;img608=8'd32;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd32;img628=8'd127;img629=8'd112;img630=8'd12;img631=8'd0;img632=8'd1;img633=8'd63;img634=8'd127;img635=8'd89;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd44;img657=8'd119;img658=8'd111;img659=8'd60;img660=8'd89;img661=8'd127;img662=8'd109;img663=8'd14;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd9;img686=8'd77;img687=8'd98;img688=8'd98;img689=8'd51;img690=8'd13;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd2;img148=8'd5;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd34;img159=8'd127;img160=8'd107;img161=8'd13;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd31;img176=8'd114;img177=8'd18;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd3;img186=8'd94;img187=8'd127;img188=8'd127;img189=8'd83;img190=8'd2;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd3;img203=8'd91;img204=8'd127;img205=8'd90;img206=8'd15;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd25;img214=8'd127;img215=8'd127;img216=8'd127;img217=8'd127;img218=8'd12;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd19;img231=8'd127;img232=8'd127;img233=8'd127;img234=8'd64;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd36;img242=8'd127;img243=8'd127;img244=8'd127;img245=8'd94;img246=8'd4;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd19;img259=8'd127;img260=8'd127;img261=8'd127;img262=8'd84;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd85;img270=8'd127;img271=8'd127;img272=8'd117;img273=8'd31;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd36;img287=8'd127;img288=8'd127;img289=8'd127;img290=8'd84;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd6;img297=8'd97;img298=8'd127;img299=8'd127;img300=8'd84;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd79;img315=8'd127;img316=8'd127;img317=8'd127;img318=8'd84;img319=8'd0;img320=8'd0;img321=8'd21;img322=8'd26;img323=8'd68;img324=8'd84;img325=8'd127;img326=8'd127;img327=8'd127;img328=8'd84;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd79;img343=8'd127;img344=8'd127;img345=8'd127;img346=8'd101;img347=8'd72;img348=8'd80;img349=8'd118;img350=8'd119;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd127;img355=8'd127;img356=8'd62;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd79;img371=8'd127;img372=8'd127;img373=8'd127;img374=8'd127;img375=8'd127;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd127;img383=8'd94;img384=8'd3;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd79;img399=8'd127;img400=8'd127;img401=8'd127;img402=8'd127;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd90;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd12;img426=8'd125;img427=8'd127;img428=8'd127;img429=8'd127;img430=8'd127;img431=8'd127;img432=8'd127;img433=8'd127;img434=8'd125;img435=8'd125;img436=8'd127;img437=8'd128;img438=8'd127;img439=8'd59;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd43;img455=8'd117;img456=8'd127;img457=8'd127;img458=8'd127;img459=8'd127;img460=8'd116;img461=8'd86;img462=8'd26;img463=8'd73;img464=8'd127;img465=8'd127;img466=8'd127;img467=8'd36;img468=8'd10;img469=8'd2;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd10;img484=8'd92;img485=8'd109;img486=8'd88;img487=8'd48;img488=8'd5;img489=8'd0;img490=8'd0;img491=8'd36;img492=8'd127;img493=8'd127;img494=8'd127;img495=8'd113;img496=8'd112;img497=8'd16;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd13;img520=8'd127;img521=8'd127;img522=8'd127;img523=8'd127;img524=8'd73;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd56;img548=8'd127;img549=8'd127;img550=8'd127;img551=8'd86;img552=8'd7;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd5;img575=8'd114;img576=8'd127;img577=8'd127;img578=8'd118;img579=8'd22;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd27;img603=8'd127;img604=8'd127;img605=8'd127;img606=8'd76;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd44;img631=8'd127;img632=8'd127;img633=8'd106;img634=8'd5;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd7;img659=8'd127;img660=8'd127;img661=8'd103;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd4;img687=8'd101;img688=8'd127;img689=8'd74;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd19;img204=8'd63;img205=8'd85;img206=8'd76;img207=8'd128;img208=8'd87;img209=8'd97;img210=8'd51;img211=8'd51;img212=8'd6;img213=8'd34;img214=8'd51;img215=8'd8;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd47;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd103;img241=8'd118;img242=8'd127;img243=8'd85;img244=8'd9;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd47;img260=8'd127;img261=8'd127;img262=8'd127;img263=8'd127;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd127;img270=8'd127;img271=8'd127;img272=8'd46;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd2;img288=8'd15;img289=8'd106;img290=8'd83;img291=8'd86;img292=8'd127;img293=8'd98;img294=8'd127;img295=8'd127;img296=8'd127;img297=8'd127;img298=8'd127;img299=8'd127;img300=8'd46;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd17;img318=8'd2;img319=8'd4;img320=8'd31;img321=8'd12;img322=8'd31;img323=8'd77;img324=8'd127;img325=8'd127;img326=8'd127;img327=8'd103;img328=8'd11;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd62;img352=8'd127;img353=8'd127;img354=8'd127;img355=8'd96;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd11;img379=8'd123;img380=8'd127;img381=8'd127;img382=8'd107;img383=8'd17;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd68;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd69;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd21;img434=8'd108;img435=8'd127;img436=8'd127;img437=8'd123;img438=8'd34;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd109;img462=8'd127;img463=8'd127;img464=8'd127;img465=8'd49;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd2;img488=8'd52;img489=8'd123;img490=8'd127;img491=8'd127;img492=8'd102;img493=8'd13;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd54;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd127;img520=8'd55;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd93;img544=8'd127;img545=8'd127;img546=8'd124;img547=8'd55;img548=8'd2;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd93;img572=8'd127;img573=8'd127;img574=8'd115;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd93;img600=8'd127;img601=8'd127;img602=8'd115;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd37;img627=8'd122;img628=8'd127;img629=8'd127;img630=8'd96;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd45;img655=8'd127;img656=8'd127;img657=8'd126;img658=8'd37;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd87;img683=8'd127;img684=8'd127;img685=8'd88;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd34;img711=8'd119;img712=8'd127;img713=8'd25;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd93;img740=8'd127;img741=8'd11;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd34;img147=8'd78;img148=8'd127;img149=8'd127;img150=8'd128;img151=8'd127;img152=8'd127;img153=8'd127;img154=8'd83;img155=8'd9;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd56;img174=8'd119;img175=8'd126;img176=8'd126;img177=8'd126;img178=8'd127;img179=8'd126;img180=8'd126;img181=8'd126;img182=8'd126;img183=8'd53;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd68;img202=8'd116;img203=8'd116;img204=8'd80;img205=8'd19;img206=8'd11;img207=8'd11;img208=8'd20;img209=8'd126;img210=8'd126;img211=8'd53;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd24;img237=8'd126;img238=8'd126;img239=8'd53;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd18;img264=8'd112;img265=8'd126;img266=8'd104;img267=8'd9;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd13;img291=8'd79;img292=8'd127;img293=8'd122;img294=8'd18;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd18;img318=8'd92;img319=8'd126;img320=8'd126;img321=8'd119;img322=8'd51;img323=8'd18;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd10;img344=8'd64;img345=8'd112;img346=8'd127;img347=8'd126;img348=8'd126;img349=8'd126;img350=8'd126;img351=8'd121;img352=8'd77;img353=8'd10;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd77;img372=8'd126;img373=8'd126;img374=8'd108;img375=8'd77;img376=8'd42;img377=8'd77;img378=8'd108;img379=8'd127;img380=8'd126;img381=8'd101;img382=8'd11;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd22;img388=8'd6;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd50;img400=8'd126;img401=8'd82;img402=8'd9;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd9;img407=8'd61;img408=8'd126;img409=8'd126;img410=8'd113;img411=8'd18;img412=8'd0;img413=8'd0;img414=8'd54;img415=8'd71;img416=8'd4;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd18;img437=8'd112;img438=8'd127;img439=8'd61;img440=8'd53;img441=8'd114;img442=8'd112;img443=8'd18;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd46;img466=8'd126;img467=8'd126;img468=8'd127;img469=8'd95;img470=8'd16;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd4;img493=8'd43;img494=8'd126;img495=8'd126;img496=8'd81;img497=8'd7;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd28;img520=8'd99;img521=8'd126;img522=8'd126;img523=8'd126;img524=8'd53;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd45;img547=8'd118;img548=8'd126;img549=8'd126;img550=8'd126;img551=8'd126;img552=8'd9;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd2;img573=8'd35;img574=8'd118;img575=8'd106;img576=8'd38;img577=8'd123;img578=8'd127;img579=8'd96;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd51;img601=8'd126;img602=8'd109;img603=8'd21;img604=8'd93;img605=8'd126;img606=8'd126;img607=8'd34;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd22;img628=8'd117;img629=8'd126;img630=8'd56;img631=8'd96;img632=8'd126;img633=8'd126;img634=8'd67;img635=8'd2;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd43;img656=8'd126;img657=8'd126;img658=8'd126;img659=8'd127;img660=8'd126;img661=8'd67;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd43;img684=8'd126;img685=8'd126;img686=8'd126;img687=8'd96;img688=8'd56;img689=8'd2;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd23;img68=8'd87;img69=8'd127;img70=8'd47;img71=8'd1;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd3;img95=8'd100;img96=8'd127;img97=8'd127;img98=8'd127;img99=8'd6;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd40;img123=8'd127;img124=8'd100;img125=8'd48;img126=8'd103;img127=8'd5;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd17;img150=8'd115;img151=8'd127;img152=8'd84;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd39;img178=8'd127;img179=8'd118;img180=8'd36;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd85;img206=8'd127;img207=8'd73;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd15;img233=8'd119;img234=8'd127;img235=8'd30;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd19;img261=8'd127;img262=8'd127;img263=8'd30;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd73;img289=8'd127;img290=8'd127;img291=8'd30;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd79;img317=8'd127;img318=8'd127;img319=8'd30;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd38;img327=8'd101;img328=8'd78;img329=8'd15;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd79;img345=8'd127;img346=8'd127;img347=8'd30;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd1;img353=8'd41;img354=8'd105;img355=8'd127;img356=8'd127;img357=8'd110;img358=8'd16;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd79;img373=8'd127;img374=8'd127;img375=8'd30;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd41;img381=8'd127;img382=8'd127;img383=8'd127;img384=8'd127;img385=8'd127;img386=8'd109;img387=8'd11;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd70;img401=8'd127;img402=8'd127;img403=8'd30;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd9;img408=8'd105;img409=8'd127;img410=8'd116;img411=8'd68;img412=8'd48;img413=8'd108;img414=8'd127;img415=8'd56;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd19;img429=8'd127;img430=8'd127;img431=8'd30;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd72;img436=8'd127;img437=8'd107;img438=8'd16;img439=8'd0;img440=8'd0;img441=8'd97;img442=8'd127;img443=8'd78;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd14;img457=8'd117;img458=8'd127;img459=8'd45;img460=8'd0;img461=8'd0;img462=8'd83;img463=8'd125;img464=8'd123;img465=8'd16;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd97;img470=8'd127;img471=8'd64;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd68;img486=8'd127;img487=8'd118;img488=8'd36;img489=8'd14;img490=8'd119;img491=8'd127;img492=8'd58;img493=8'd0;img494=8'd0;img495=8'd7;img496=8'd51;img497=8'd120;img498=8'd94;img499=8'd5;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd17;img514=8'd115;img515=8'd127;img516=8'd119;img517=8'd112;img518=8'd127;img519=8'd127;img520=8'd0;img521=8'd0;img522=8'd27;img523=8'd88;img524=8'd127;img525=8'd127;img526=8'd64;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd28;img543=8'd116;img544=8'd127;img545=8'd127;img546=8'd127;img547=8'd127;img548=8'd107;img549=8'd83;img550=8'd120;img551=8'd127;img552=8'd127;img553=8'd72;img554=8'd4;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd56;img572=8'd117;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd127;img579=8'd116;img580=8'd58;img581=8'd3;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd5;img601=8'd58;img602=8'd66;img603=8'd124;img604=8'd127;img605=8'd121;img606=8'd66;img607=8'd25;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd60;img129=8'd127;img130=8'd108;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd59;img157=8'd127;img158=8'd107;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd0;img183=8'd0;img184=8'd59;img185=8'd127;img186=8'd107;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd0;img210=8'd0;img211=8'd5;img212=8'd69;img213=8'd127;img214=8'd107;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd0;img237=8'd0;img238=8'd0;img239=8'd67;img240=8'd127;img241=8'd127;img242=8'd107;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd127;img268=8'd127;img269=8'd127;img270=8'd47;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd84;img295=8'd128;img296=8'd127;img297=8'd52;img298=8'd2;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd22;img322=8'd107;img323=8'd127;img324=8'd108;img325=8'd27;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd22;img349=8'd100;img350=8'd127;img351=8'd127;img352=8'd68;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd40;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd68;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd10;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd122;img408=8'd53;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd6;img432=8'd86;img433=8'd127;img434=8'd127;img435=8'd112;img436=8'd32;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd40;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd68;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd10;img488=8'd120;img489=8'd127;img490=8'd127;img491=8'd100;img492=8'd5;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd48;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd61;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd108;img544=8'd127;img545=8'd127;img546=8'd127;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd67;img571=8'd124;img572=8'd127;img573=8'd127;img574=8'd119;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd78;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd29;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd78;img627=8'd127;img628=8'd127;img629=8'd127;img630=8'd29;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd18;img655=8'd37;img656=8'd96;img657=8'd29;img658=8'd7;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd11;img153=8'd58;img154=8'd98;img155=8'd127;img156=8'd127;img157=8'd127;img158=8'd78;img159=8'd9;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd33;img180=8'd102;img181=8'd127;img182=8'd127;img183=8'd126;img184=8'd124;img185=8'd127;img186=8'd127;img187=8'd80;img188=8'd1;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd4;img206=8'd69;img207=8'd125;img208=8'd127;img209=8'd121;img210=8'd74;img211=8'd34;img212=8'd21;img213=8'd59;img214=8'd123;img215=8'd127;img216=8'd10;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd55;img234=8'd127;img235=8'd121;img236=8'd79;img237=8'd15;img238=8'd0;img239=8'd0;img240=8'd1;img241=8'd58;img242=8'd125;img243=8'd124;img244=8'd9;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd11;img262=8'd73;img263=8'd18;img264=8'd0;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd23;img269=8'd127;img270=8'd127;img271=8'd53;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd0;img293=8'd3;img294=8'd56;img295=8'd77;img296=8'd120;img297=8'd127;img298=8'd110;img299=8'd4;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd42;img322=8'd127;img323=8'd127;img324=8'd127;img325=8'd115;img326=8'd24;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd74;img348=8'd120;img349=8'd124;img350=8'd127;img351=8'd127;img352=8'd127;img353=8'd125;img354=8'd50;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd120;img376=8'd127;img377=8'd127;img378=8'd126;img379=8'd91;img380=8'd127;img381=8'd127;img382=8'd124;img383=8'd48;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd2;img404=8'd22;img405=8'd2;img406=8'd2;img407=8'd1;img408=8'd25;img409=8'd92;img410=8'd127;img411=8'd126;img412=8'd39;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd7;img438=8'd114;img439=8'd127;img440=8'd61;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd63;img467=8'd127;img468=8'd110;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd65;img495=8'd127;img496=8'd107;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd54;img512=8'd47;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd0;img521=8'd0;img522=8'd112;img523=8'd127;img524=8'd60;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd16;img539=8'd118;img540=8'd84;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd1;img549=8'd60;img550=8'd125;img551=8'd127;img552=8'd35;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd33;img567=8'd127;img568=8'd89;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd24;img577=8'd127;img578=8'd127;img579=8'd83;img580=8'd3;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd16;img595=8'd118;img596=8'd89;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd9;img603=8'd79;img604=8'd122;img605=8'd127;img606=8'd102;img607=8'd3;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd110;img624=8'd118;img625=8'd69;img626=8'd45;img627=8'd45;img628=8'd46;img629=8'd75;img630=8'd108;img631=8'd127;img632=8'd124;img633=8'd82;img634=8'd10;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd81;img652=8'd127;img653=8'd127;img654=8'd127;img655=8'd127;img656=8'd127;img657=8'd127;img658=8'd118;img659=8'd73;img660=8'd12;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd13;img680=8'd62;img681=8'd83;img682=8'd127;img683=8'd99;img684=8'd77;img685=8'd67;img686=8'd16;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd7;img72=8'd71;img73=8'd112;img74=8'd40;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd93;img100=8'd127;img101=8'd127;img102=8'd59;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd50;img127=8'd127;img128=8'd86;img129=8'd58;img130=8'd18;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd26;img154=8'd124;img155=8'd122;img156=8'd20;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd16;img181=8'd110;img182=8'd127;img183=8'd23;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd3;img208=8'd60;img209=8'd127;img210=8'd86;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd52;img236=8'd127;img237=8'd106;img238=8'd5;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd10;img263=8'd98;img264=8'd114;img265=8'd22;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd75;img291=8'd127;img292=8'd87;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd97;img319=8'd127;img320=8'd50;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd12;img346=8'd128;img347=8'd87;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd25;img353=8'd49;img354=8'd30;img355=8'd7;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd90;img374=8'd127;img375=8'd68;img376=8'd0;img377=8'd0;img378=8'd27;img379=8'd108;img380=8'd124;img381=8'd127;img382=8'd127;img383=8'd93;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd98;img402=8'd127;img403=8'd68;img404=8'd0;img405=8'd44;img406=8'd118;img407=8'd127;img408=8'd108;img409=8'd54;img410=8'd86;img411=8'd127;img412=8'd34;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd98;img430=8'd127;img431=8'd68;img432=8'd44;img433=8'd126;img434=8'd127;img435=8'd77;img436=8'd13;img437=8'd0;img438=8'd68;img439=8'd127;img440=8'd87;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd98;img458=8'd127;img459=8'd75;img460=8'd118;img461=8'd119;img462=8'd59;img463=8'd0;img464=8'd0;img465=8'd0;img466=8'd68;img467=8'd127;img468=8'd49;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd50;img486=8'd128;img487=8'd127;img488=8'd127;img489=8'd77;img490=8'd0;img491=8'd0;img492=8'd0;img493=8'd0;img494=8'd69;img495=8'd127;img496=8'd12;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd8;img514=8'd104;img515=8'd127;img516=8'd127;img517=8'd62;img518=8'd0;img519=8'd7;img520=8'd10;img521=8'd10;img522=8'd92;img523=8'd123;img524=8'd27;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd64;img543=8'd127;img544=8'd127;img545=8'd121;img546=8'd88;img547=8'd112;img548=8'd127;img549=8'd127;img550=8'd127;img551=8'd63;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd3;img571=8'd55;img572=8'd121;img573=8'd127;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd108;img579=8'd3;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd21;img601=8'd82;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd111;img606=8'd47;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd0;img182=8'd3;img183=8'd58;img184=8'd122;img185=8'd112;img186=8'd123;img187=8'd30;img188=8'd0;img189=8'd16;img190=8'd61;img191=8'd1;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd0;img209=8'd1;img210=8'd75;img211=8'd96;img212=8'd48;img213=8'd4;img214=8'd79;img215=8'd13;img216=8'd9;img217=8'd110;img218=8'd114;img219=8'd11;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd0;img236=8'd7;img237=8'd87;img238=8'd75;img239=8'd28;img240=8'd0;img241=8'd0;img242=8'd31;img243=8'd3;img244=8'd99;img245=8'd114;img246=8'd22;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd0;img264=8'd43;img265=8'd100;img266=8'd13;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd33;img272=8'd102;img273=8'd38;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd63;img293=8'd69;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd22;img299=8'd122;img300=8'd115;img301=8'd23;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd70;img320=8'd101;img321=8'd3;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd75;img327=8'd126;img328=8'd42;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd44;img347=8'd114;img348=8'd5;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd9;img353=8'd76;img354=8'd127;img355=8'd70;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd2;img374=8'd113;img375=8'd48;img376=8'd0;img377=8'd0;img378=8'd1;img379=8'd34;img380=8'd97;img381=8'd112;img382=8'd55;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd25;img402=8'd115;img403=8'd10;img404=8'd14;img405=8'd30;img406=8'd76;img407=8'd128;img408=8'd125;img409=8'd36;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd21;img430=8'd125;img431=8'd103;img432=8'd127;img433=8'd111;img434=8'd103;img435=8'd123;img436=8'd101;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd53;img459=8'd98;img460=8'd62;img461=8'd8;img462=8'd68;img463=8'd123;img464=8'd71;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd55;img490=8'd127;img491=8'd99;img492=8'd3;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd15;img517=8'd125;img518=8'd119;img519=8'd13;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd2;img544=8'd110;img545=8'd105;img546=8'd12;img547=8'd0;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd56;img572=8'd122;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd32;img599=8'd122;img600=8'd62;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd47;img626=8'd117;img627=8'd82;img628=8'd2;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd106;img654=8'd111;img655=8'd5;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd106;img682=8'd63;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd12;img709=8'd45;img710=8'd1;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd55;img150=8'd63;img151=8'd63;img152=8'd63;img153=8'd79;img154=8'd79;img155=8'd63;img156=8'd19;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd79;img177=8'd127;img178=8'd127;img179=8'd127;img180=8'd127;img181=8'd128;img182=8'd127;img183=8'd127;img184=8'd126;img185=8'd42;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd86;img205=8'd127;img206=8'd127;img207=8'd127;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd124;img214=8'd72;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd4;img233=8'd52;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd111;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd5;img262=8'd13;img263=8'd67;img264=8'd92;img265=8'd127;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd127;img270=8'd111;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd92;img292=8'd116;img293=8'd127;img294=8'd127;img295=8'd127;img296=8'd127;img297=8'd127;img298=8'd111;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd59;img319=8'd124;img320=8'd127;img321=8'd127;img322=8'd127;img323=8'd127;img324=8'd127;img325=8'd127;img326=8'd56;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd108;img347=8'd127;img348=8'd127;img349=8'd127;img350=8'd127;img351=8'd127;img352=8'd127;img353=8'd127;img354=8'd66;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd44;img375=8'd121;img376=8'd127;img377=8'd127;img378=8'd127;img379=8'd127;img380=8'd127;img381=8'd127;img382=8'd111;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd45;img404=8'd121;img405=8'd127;img406=8'd103;img407=8'd118;img408=8'd127;img409=8'd127;img410=8'd115;img411=8'd13;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd26;img433=8'd33;img434=8'd9;img435=8'd77;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd64;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd27;img464=8'd127;img465=8'd127;img466=8'd127;img467=8'd114;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd0;img491=8'd39;img492=8'd127;img493=8'd127;img494=8'd127;img495=8'd69;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd20;img519=8'd116;img520=8'd127;img521=8'd127;img522=8'd127;img523=8'd49;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd9;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd5;img546=8'd76;img547=8'd127;img548=8'd127;img549=8'd127;img550=8'd117;img551=8'd18;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd71;img569=8'd104;img570=8'd79;img571=8'd25;img572=8'd66;img573=8'd91;img574=8'd127;img575=8'd127;img576=8'd127;img577=8'd127;img578=8'd104;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd32;img596=8'd122;img597=8'd127;img598=8'd127;img599=8'd127;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd127;img605=8'd126;img606=8'd42;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd53;img624=8'd127;img625=8'd127;img626=8'd127;img627=8'd127;img628=8'd127;img629=8'd127;img630=8'd127;img631=8'd127;img632=8'd123;img633=8'd68;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd25;img652=8'd118;img653=8'd127;img654=8'd127;img655=8'd127;img656=8'd127;img657=8'd127;img658=8'd125;img659=8'd111;img660=8'd18;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd55;img682=8'd118;img683=8'd127;img684=8'd127;img685=8'd111;img686=8'd16;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd46;img124=8'd127;img125=8'd127;img126=8'd127;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd95;img152=8'd126;img153=8'd126;img154=8'd126;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd95;img180=8'd126;img181=8'd126;img182=8'd126;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd95;img208=8'd126;img209=8'd126;img210=8'd126;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd95;img236=8'd126;img237=8'd126;img238=8'd126;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd96;img264=8'd127;img265=8'd127;img266=8'd127;img267=8'd98;img268=8'd12;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd95;img292=8'd126;img293=8'd126;img294=8'd126;img295=8'd127;img296=8'd31;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd95;img320=8'd126;img321=8'd126;img322=8'd126;img323=8'd127;img324=8'd71;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd26;img348=8'd126;img349=8'd126;img350=8'd126;img351=8'd127;img352=8'd110;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd16;img376=8'd126;img377=8'd126;img378=8'd126;img379=8'd127;img380=8'd110;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd6;img404=8'd87;img405=8'd127;img406=8'd127;img407=8'd128;img408=8'd111;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd16;img432=8'd126;img433=8'd126;img434=8'd126;img435=8'd127;img436=8'd110;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd16;img460=8'd126;img461=8'd126;img462=8'd126;img463=8'd127;img464=8'd110;img465=8'd0;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd16;img488=8'd126;img489=8'd126;img490=8'd126;img491=8'd127;img492=8'd110;img493=8'd0;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd16;img516=8'd126;img517=8'd126;img518=8'd126;img519=8'd127;img520=8'd110;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd10;img544=8'd103;img545=8'd127;img546=8'd127;img547=8'd128;img548=8'd127;img549=8'd63;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd16;img573=8'd115;img574=8'd126;img575=8'd127;img576=8'd126;img577=8'd63;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd111;img602=8'd126;img603=8'd127;img604=8'd126;img605=8'd94;img606=8'd48;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd91;img630=8'd106;img631=8'd127;img632=8'd126;img633=8'd126;img634=8'd94;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd12;img658=8'd18;img659=8'd77;img660=8'd126;img661=8'd126;img662=8'd45;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd19;img159=8'd127;img160=8'd128;img161=8'd127;img162=8'd36;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd0;img181=8'd32;img182=8'd32;img183=8'd0;img184=8'd0;img185=8'd32;img186=8'd91;img187=8'd126;img188=8'd127;img189=8'd126;img190=8'd36;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd0;img208=8'd91;img209=8'd121;img210=8'd108;img211=8'd0;img212=8'd8;img213=8'd111;img214=8'd126;img215=8'd126;img216=8'd119;img217=8'd87;img218=8'd10;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd11;img235=8'd72;img236=8'd127;img237=8'd105;img238=8'd46;img239=8'd1;img240=8'd96;img241=8'd126;img242=8'd126;img243=8'd126;img244=8'd72;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd47;img262=8'd106;img263=8'd126;img264=8'd103;img265=8'd10;img266=8'd0;img267=8'd72;img268=8'd127;img269=8'd126;img270=8'd126;img271=8'd54;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd16;img289=8'd114;img290=8'd126;img291=8'd126;img292=8'd10;img293=8'd0;img294=8'd16;img295=8'd119;img296=8'd127;img297=8'd126;img298=8'd110;img299=8'd8;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd3;img315=8'd19;img316=8'd106;img317=8'd126;img318=8'd123;img319=8'd66;img320=8'd0;img321=8'd6;img322=8'd75;img323=8'd126;img324=8'd127;img325=8'd126;img326=8'd98;img327=8'd0;img328=8'd0;img329=8'd11;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd19;img343=8'd126;img344=8'd126;img345=8'd126;img346=8'd66;img347=8'd0;img348=8'd0;img349=8'd37;img350=8'd126;img351=8'd126;img352=8'd127;img353=8'd126;img354=8'd36;img355=8'd0;img356=8'd73;img357=8'd103;img358=8'd21;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd91;img371=8'd127;img372=8'd127;img373=8'd127;img374=8'd36;img375=8'd0;img376=8'd0;img377=8'd37;img378=8'd127;img379=8'd127;img380=8'd128;img381=8'd106;img382=8'd55;img383=8'd96;img384=8'd128;img385=8'd127;img386=8'd36;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd32;img398=8'd121;img399=8'd126;img400=8'd126;img401=8'd126;img402=8'd62;img403=8'd37;img404=8'd21;img405=8'd58;img406=8'd126;img407=8'd126;img408=8'd127;img409=8'd126;img410=8'd126;img411=8'd126;img412=8'd127;img413=8'd116;img414=8'd26;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd37;img426=8'd126;img427=8'd126;img428=8'd126;img429=8'd126;img430=8'd126;img431=8'd126;img432=8'd111;img433=8'd121;img434=8'd126;img435=8'd126;img436=8'd127;img437=8'd126;img438=8'd126;img439=8'd126;img440=8'd119;img441=8'd77;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd37;img454=8'd126;img455=8'd126;img456=8'd126;img457=8'd126;img458=8'd126;img459=8'd126;img460=8'd127;img461=8'd126;img462=8'd126;img463=8'd126;img464=8'd127;img465=8'd126;img466=8'd126;img467=8'd126;img468=8'd72;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd21;img482=8'd80;img483=8'd127;img484=8'd127;img485=8'd127;img486=8'd127;img487=8'd127;img488=8'd128;img489=8'd127;img490=8'd127;img491=8'd127;img492=8'd128;img493=8'd127;img494=8'd119;img495=8'd72;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd3;img511=8'd60;img512=8'd105;img513=8'd95;img514=8'd116;img515=8'd126;img516=8'd127;img517=8'd126;img518=8'd126;img519=8'd126;img520=8'd111;img521=8'd69;img522=8'd15;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd16;img541=8'd5;img542=8'd26;img543=8'd77;img544=8'd127;img545=8'd126;img546=8'd126;img547=8'd126;img548=8'd80;img549=8'd3;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd127;img573=8'd126;img574=8'd126;img575=8'd126;img576=8'd127;img577=8'd60;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd96;img601=8'd127;img602=8'd127;img603=8'd127;img604=8'd128;img605=8'd127;img606=8'd67;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd39;img629=8'd121;img630=8'd126;img631=8'd126;img632=8'd127;img633=8'd126;img634=8'd87;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd52;img658=8'd111;img659=8'd126;img660=8'd127;img661=8'd110;img662=8'd31;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd8;img687=8'd95;img688=8'd54;img689=8'd8;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd11;img150=8'd123;img151=8'd43;img152=8'd3;img153=8'd6;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd40;img179=8'd120;img180=8'd89;img181=8'd102;img182=8'd0;img183=8'd0;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd92;img208=8'd126;img209=8'd126;img210=8'd0;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd0;img235=8'd92;img236=8'd126;img237=8'd126;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd0;img262=8'd0;img263=8'd66;img264=8'd126;img265=8'd126;img266=8'd53;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd16;img292=8'd115;img293=8'd127;img294=8'd122;img295=8'd25;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd67;img321=8'd126;img322=8'd127;img323=8'd57;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd34;img349=8'd108;img350=8'd127;img351=8'd110;img352=8'd10;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd0;img373=8'd0;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd11;img378=8'd127;img379=8'd126;img380=8'd56;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd0;img401=8'd0;img402=8'd0;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd127;img407=8'd126;img408=8'd92;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd0;img430=8'd0;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd128;img435=8'd127;img436=8'd92;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd80;img463=8'd126;img464=8'd98;img465=8'd5;img466=8'd0;img467=8'd0;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd0;img488=8'd0;img489=8'd0;img490=8'd9;img491=8'd114;img492=8'd126;img493=8'd23;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd0;img516=8'd0;img517=8'd0;img518=8'd0;img519=8'd81;img520=8'd126;img521=8'd23;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd29;img548=8'd126;img549=8'd75;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd24;img576=8'd127;img577=8'd81;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd24;img604=8'd126;img605=8'd80;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd24;img632=8'd126;img633=8'd80;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd24;img660=8'd126;img661=8'd118;img662=8'd10;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd3;img688=8'd69;img689=8'd58;img690=8'd1;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd14;img176=8'd68;img177=8'd29;img178=8'd9;img179=8'd9;img180=8'd9;img181=8'd9;img182=8'd9;img183=8'd19;img184=8'd68;img185=8'd23;img186=8'd2;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd127;img204=8'd127;img205=8'd127;img206=8'd127;img207=8'd127;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd127;img214=8'd21;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd128;img232=8'd127;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd127;img238=8'd127;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd21;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd37;img260=8'd91;img261=8'd79;img262=8'd33;img263=8'd81;img264=8'd106;img265=8'd127;img266=8'd127;img267=8'd127;img268=8'd127;img269=8'd116;img270=8'd15;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd0;img290=8'd0;img291=8'd0;img292=8'd29;img293=8'd124;img294=8'd127;img295=8'd127;img296=8'd117;img297=8'd30;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd0;img317=8'd0;img318=8'd0;img319=8'd0;img320=8'd6;img321=8'd122;img322=8'd127;img323=8'd127;img324=8'd124;img325=8'd26;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd0;img345=8'd0;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd94;img350=8'd127;img351=8'd127;img352=8'd97;img353=8'd2;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd2;img373=8'd12;img374=8'd57;img375=8'd71;img376=8'd71;img377=8'd125;img378=8'd127;img379=8'd127;img380=8'd47;img381=8'd12;img382=8'd12;img383=8'd12;img384=8'd12;img385=8'd12;img386=8'd12;img387=8'd12;img388=8'd12;img389=8'd12;img390=8'd7;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd15;img401=8'd120;img402=8'd127;img403=8'd127;img404=8'd127;img405=8'd127;img406=8'd127;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd127;img413=8'd127;img414=8'd127;img415=8'd127;img416=8'd127;img417=8'd119;img418=8'd84;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd0;img429=8'd26;img430=8'd55;img431=8'd108;img432=8'd127;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd127;img440=8'd127;img441=8'd127;img442=8'd108;img443=8'd97;img444=8'd78;img445=8'd23;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd0;img456=8'd0;img457=8'd0;img458=8'd0;img459=8'd45;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd121;img464=8'd115;img465=8'd97;img466=8'd88;img467=8'd35;img468=8'd30;img469=8'd30;img470=8'd11;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd0;img484=8'd0;img485=8'd0;img486=8'd0;img487=8'd45;img488=8'd127;img489=8'd127;img490=8'd127;img491=8'd84;img492=8'd15;img493=8'd5;img494=8'd0;img495=8'd0;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd0;img515=8'd45;img516=8'd127;img517=8'd127;img518=8'd127;img519=8'd47;img520=8'd0;img521=8'd0;img522=8'd0;img523=8'd0;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd45;img544=8'd127;img545=8'd127;img546=8'd115;img547=8'd1;img548=8'd0;img549=8'd0;img550=8'd0;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd45;img572=8'd127;img573=8'd127;img574=8'd122;img575=8'd28;img576=8'd0;img577=8'd0;img578=8'd0;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd45;img600=8'd127;img601=8'd127;img602=8'd127;img603=8'd47;img604=8'd0;img605=8'd0;img606=8'd0;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd45;img628=8'd127;img629=8'd127;img630=8'd127;img631=8'd47;img632=8'd0;img633=8'd0;img634=8'd0;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd45;img656=8'd127;img657=8'd127;img658=8'd117;img659=8'd10;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd45;img684=8'd127;img685=8'd127;img686=8'd115;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd3;img712=8'd61;img713=8'd68;img714=8'd34;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd11;img100=8'd79;img101=8'd121;img102=8'd124;img103=8'd65;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd2;img126=8'd44;img127=8'd121;img128=8'd121;img129=8'd99;img130=8'd111;img131=8'd127;img132=8'd76;img133=8'd2;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd10;img153=8'd84;img154=8'd127;img155=8'd122;img156=8'd21;img157=8'd0;img158=8'd8;img159=8'd89;img160=8'd127;img161=8'd55;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd0;img178=8'd0;img179=8'd0;img180=8'd73;img181=8'd127;img182=8'd104;img183=8'd20;img184=8'd0;img185=8'd0;img186=8'd0;img187=8'd26;img188=8'd118;img189=8'd60;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd0;img205=8'd0;img206=8'd0;img207=8'd36;img208=8'd122;img209=8'd120;img210=8'd11;img211=8'd0;img212=8'd0;img213=8'd0;img214=8'd0;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd0;img232=8'd0;img233=8'd0;img234=8'd11;img235=8'd105;img236=8'd122;img237=8'd36;img238=8'd0;img239=8'd0;img240=8'd0;img241=8'd0;img242=8'd0;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd0;img259=8'd0;img260=8'd0;img261=8'd10;img262=8'd105;img263=8'd127;img264=8'd73;img265=8'd0;img266=8'd0;img267=8'd0;img268=8'd0;img269=8'd0;img270=8'd0;img271=8'd0;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd0;img287=8'd0;img288=8'd0;img289=8'd68;img290=8'd127;img291=8'd113;img292=8'd9;img293=8'd0;img294=8'd0;img295=8'd0;img296=8'd0;img297=8'd0;img298=8'd0;img299=8'd0;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd0;img315=8'd0;img316=8'd11;img317=8'd119;img318=8'd127;img319=8'd45;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd0;img325=8'd0;img326=8'd0;img327=8'd0;img328=8'd0;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd0;img343=8'd0;img344=8'd55;img345=8'd127;img346=8'd101;img347=8'd3;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd0;img352=8'd0;img353=8'd0;img354=8'd0;img355=8'd0;img356=8'd0;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd0;img371=8'd0;img372=8'd68;img373=8'd127;img374=8'd91;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd0;img379=8'd0;img380=8'd0;img381=8'd0;img382=8'd0;img383=8'd0;img384=8'd0;img385=8'd0;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd0;img399=8'd0;img400=8'd58;img401=8'd127;img402=8'd65;img403=8'd0;img404=8'd0;img405=8'd0;img406=8'd0;img407=8'd0;img408=8'd0;img409=8'd0;img410=8'd0;img411=8'd0;img412=8'd0;img413=8'd0;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd0;img427=8'd0;img428=8'd77;img429=8'd127;img430=8'd46;img431=8'd0;img432=8'd0;img433=8'd0;img434=8'd0;img435=8'd0;img436=8'd0;img437=8'd0;img438=8'd0;img439=8'd0;img440=8'd0;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd0;img455=8'd14;img456=8'd119;img457=8'd127;img458=8'd65;img459=8'd0;img460=8'd0;img461=8'd0;img462=8'd0;img463=8'd6;img464=8'd10;img465=8'd10;img466=8'd10;img467=8'd6;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd14;img484=8'd119;img485=8'd127;img486=8'd91;img487=8'd0;img488=8'd0;img489=8'd20;img490=8'd62;img491=8'd114;img492=8'd127;img493=8'd127;img494=8'd127;img495=8'd114;img496=8'd33;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd71;img513=8'd127;img514=8'd101;img515=8'd3;img516=8'd77;img517=8'd127;img518=8'd127;img519=8'd128;img520=8'd93;img521=8'd96;img522=8'd127;img523=8'd127;img524=8'd101;img525=8'd3;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd45;img541=8'd127;img542=8'd127;img543=8'd119;img544=8'd125;img545=8'd112;img546=8'd54;img547=8'd9;img548=8'd1;img549=8'd2;img550=8'd102;img551=8'd127;img552=8'd127;img553=8'd9;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd2;img569=8'd73;img570=8'd127;img571=8'd127;img572=8'd127;img573=8'd63;img574=8'd0;img575=8'd0;img576=8'd4;img577=8'd25;img578=8'd113;img579=8'd127;img580=8'd73;img581=8'd2;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd10;img598=8'd104;img599=8'd127;img600=8'd127;img601=8'd125;img602=8'd100;img603=8'd100;img604=8'd106;img605=8'd127;img606=8'd126;img607=8'd85;img608=8'd10;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd11;img627=8'd62;img628=8'd88;img629=8'd127;img630=8'd127;img631=8'd127;img632=8'd127;img633=8'd104;img634=8'd43;img635=8'd0;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd0;img661=8'd0;img662=8'd0;img663=8'd0;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd0;img689=8'd0;img690=8'd0;img691=8'd0;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd0;img717=8'd0;img718=8'd0;img719=8'd0;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
@(negedge clk)#(10/4) img0=8'd0;img1=8'd0;img2=8'd0;img3=8'd0;img4=8'd0;img5=8'd0;img6=8'd0;img7=8'd0;img8=8'd0;img9=8'd0;img10=8'd0;img11=8'd0;img12=8'd0;img13=8'd0;img14=8'd0;img15=8'd0;img16=8'd0;img17=8'd0;img18=8'd0;img19=8'd0;img20=8'd0;img21=8'd0;img22=8'd0;img23=8'd0;img24=8'd0;img25=8'd0;img26=8'd0;img27=8'd0;img28=8'd0;img29=8'd0;img30=8'd0;img31=8'd0;img32=8'd0;img33=8'd0;img34=8'd0;img35=8'd0;img36=8'd0;img37=8'd0;img38=8'd0;img39=8'd0;img40=8'd0;img41=8'd0;img42=8'd0;img43=8'd0;img44=8'd0;img45=8'd0;img46=8'd0;img47=8'd0;img48=8'd0;img49=8'd0;img50=8'd0;img51=8'd0;img52=8'd0;img53=8'd0;img54=8'd0;img55=8'd0;img56=8'd0;img57=8'd0;img58=8'd0;img59=8'd0;img60=8'd0;img61=8'd0;img62=8'd0;img63=8'd0;img64=8'd0;img65=8'd0;img66=8'd0;img67=8'd0;img68=8'd0;img69=8'd0;img70=8'd0;img71=8'd0;img72=8'd0;img73=8'd0;img74=8'd0;img75=8'd0;img76=8'd0;img77=8'd0;img78=8'd0;img79=8'd0;img80=8'd0;img81=8'd0;img82=8'd0;img83=8'd0;img84=8'd0;img85=8'd0;img86=8'd0;img87=8'd0;img88=8'd0;img89=8'd0;img90=8'd0;img91=8'd0;img92=8'd0;img93=8'd0;img94=8'd0;img95=8'd0;img96=8'd0;img97=8'd0;img98=8'd0;img99=8'd0;img100=8'd0;img101=8'd0;img102=8'd0;img103=8'd0;img104=8'd0;img105=8'd0;img106=8'd0;img107=8'd0;img108=8'd0;img109=8'd0;img110=8'd0;img111=8'd0;img112=8'd0;img113=8'd0;img114=8'd0;img115=8'd0;img116=8'd0;img117=8'd0;img118=8'd0;img119=8'd0;img120=8'd0;img121=8'd0;img122=8'd0;img123=8'd0;img124=8'd0;img125=8'd0;img126=8'd0;img127=8'd0;img128=8'd0;img129=8'd0;img130=8'd0;img131=8'd0;img132=8'd0;img133=8'd0;img134=8'd0;img135=8'd0;img136=8'd0;img137=8'd0;img138=8'd0;img139=8'd0;img140=8'd0;img141=8'd0;img142=8'd0;img143=8'd0;img144=8'd0;img145=8'd0;img146=8'd0;img147=8'd0;img148=8'd0;img149=8'd0;img150=8'd0;img151=8'd0;img152=8'd0;img153=8'd0;img154=8'd0;img155=8'd0;img156=8'd0;img157=8'd0;img158=8'd0;img159=8'd0;img160=8'd0;img161=8'd0;img162=8'd0;img163=8'd0;img164=8'd0;img165=8'd0;img166=8'd0;img167=8'd0;img168=8'd0;img169=8'd0;img170=8'd0;img171=8'd0;img172=8'd0;img173=8'd0;img174=8'd0;img175=8'd0;img176=8'd0;img177=8'd1;img178=8'd19;img179=8'd61;img180=8'd123;img181=8'd128;img182=8'd128;img183=8'd123;img184=8'd61;img185=8'd4;img186=8'd0;img187=8'd0;img188=8'd0;img189=8'd0;img190=8'd0;img191=8'd0;img192=8'd0;img193=8'd0;img194=8'd0;img195=8'd0;img196=8'd0;img197=8'd0;img198=8'd0;img199=8'd0;img200=8'd0;img201=8'd0;img202=8'd0;img203=8'd0;img204=8'd29;img205=8'd88;img206=8'd127;img207=8'd127;img208=8'd127;img209=8'd127;img210=8'd127;img211=8'd127;img212=8'd127;img213=8'd78;img214=8'd2;img215=8'd0;img216=8'd0;img217=8'd0;img218=8'd0;img219=8'd0;img220=8'd0;img221=8'd0;img222=8'd0;img223=8'd0;img224=8'd0;img225=8'd0;img226=8'd0;img227=8'd0;img228=8'd0;img229=8'd0;img230=8'd0;img231=8'd1;img232=8'd96;img233=8'd127;img234=8'd127;img235=8'd127;img236=8'd127;img237=8'd125;img238=8'd124;img239=8'd127;img240=8'd127;img241=8'd127;img242=8'd53;img243=8'd0;img244=8'd0;img245=8'd0;img246=8'd0;img247=8'd0;img248=8'd0;img249=8'd0;img250=8'd0;img251=8'd0;img252=8'd0;img253=8'd0;img254=8'd0;img255=8'd0;img256=8'd0;img257=8'd0;img258=8'd1;img259=8'd63;img260=8'd127;img261=8'd127;img262=8'd123;img263=8'd105;img264=8'd56;img265=8'd19;img266=8'd0;img267=8'd78;img268=8'd127;img269=8'd127;img270=8'd94;img271=8'd7;img272=8'd0;img273=8'd0;img274=8'd0;img275=8'd0;img276=8'd0;img277=8'd0;img278=8'd0;img279=8'd0;img280=8'd0;img281=8'd0;img282=8'd0;img283=8'd0;img284=8'd0;img285=8'd0;img286=8'd3;img287=8'd127;img288=8'd127;img289=8'd125;img290=8'd70;img291=8'd0;img292=8'd0;img293=8'd0;img294=8'd0;img295=8'd8;img296=8'd113;img297=8'd127;img298=8'd127;img299=8'd58;img300=8'd0;img301=8'd0;img302=8'd0;img303=8'd0;img304=8'd0;img305=8'd0;img306=8'd0;img307=8'd0;img308=8'd0;img309=8'd0;img310=8'd0;img311=8'd0;img312=8'd0;img313=8'd0;img314=8'd3;img315=8'd127;img316=8'd127;img317=8'd71;img318=8'd0;img319=8'd0;img320=8'd0;img321=8'd0;img322=8'd0;img323=8'd0;img324=8'd38;img325=8'd127;img326=8'd127;img327=8'd110;img328=8'd13;img329=8'd0;img330=8'd0;img331=8'd0;img332=8'd0;img333=8'd0;img334=8'd0;img335=8'd0;img336=8'd0;img337=8'd0;img338=8'd0;img339=8'd0;img340=8'd0;img341=8'd0;img342=8'd37;img343=8'd127;img344=8'd119;img345=8'd11;img346=8'd0;img347=8'd0;img348=8'd0;img349=8'd0;img350=8'd0;img351=8'd7;img352=8'd111;img353=8'd127;img354=8'd127;img355=8'd127;img356=8'd75;img357=8'd0;img358=8'd0;img359=8'd0;img360=8'd0;img361=8'd0;img362=8'd0;img363=8'd0;img364=8'd0;img365=8'd0;img366=8'd0;img367=8'd0;img368=8'd0;img369=8'd0;img370=8'd57;img371=8'd127;img372=8'd118;img373=8'd11;img374=8'd0;img375=8'd0;img376=8'd0;img377=8'd0;img378=8'd16;img379=8'd97;img380=8'd127;img381=8'd127;img382=8'd127;img383=8'd127;img384=8'd115;img385=8'd2;img386=8'd0;img387=8'd0;img388=8'd0;img389=8'd0;img390=8'd0;img391=8'd0;img392=8'd0;img393=8'd0;img394=8'd0;img395=8'd0;img396=8'd0;img397=8'd0;img398=8'd31;img399=8'd127;img400=8'd127;img401=8'd63;img402=8'd0;img403=8'd0;img404=8'd1;img405=8'd20;img406=8'd86;img407=8'd127;img408=8'd127;img409=8'd127;img410=8'd127;img411=8'd127;img412=8'd80;img413=8'd1;img414=8'd0;img415=8'd0;img416=8'd0;img417=8'd0;img418=8'd0;img419=8'd0;img420=8'd0;img421=8'd0;img422=8'd0;img423=8'd0;img424=8'd0;img425=8'd0;img426=8'd3;img427=8'd127;img428=8'd127;img429=8'd106;img430=8'd48;img431=8'd28;img432=8'd80;img433=8'd127;img434=8'd127;img435=8'd127;img436=8'd127;img437=8'd127;img438=8'd127;img439=8'd120;img440=8'd37;img441=8'd0;img442=8'd0;img443=8'd0;img444=8'd0;img445=8'd0;img446=8'd0;img447=8'd0;img448=8'd0;img449=8'd0;img450=8'd0;img451=8'd0;img452=8'd0;img453=8'd0;img454=8'd1;img455=8'd67;img456=8'd127;img457=8'd127;img458=8'd127;img459=8'd127;img460=8'd127;img461=8'd127;img462=8'd127;img463=8'd127;img464=8'd107;img465=8'd127;img466=8'd127;img467=8'd94;img468=8'd0;img469=8'd0;img470=8'd0;img471=8'd0;img472=8'd0;img473=8'd0;img474=8'd0;img475=8'd0;img476=8'd0;img477=8'd0;img478=8'd0;img479=8'd0;img480=8'd0;img481=8'd0;img482=8'd0;img483=8'd2;img484=8'd49;img485=8'd87;img486=8'd123;img487=8'd127;img488=8'd126;img489=8'd116;img490=8'd96;img491=8'd11;img492=8'd33;img493=8'd127;img494=8'd127;img495=8'd44;img496=8'd0;img497=8'd0;img498=8'd0;img499=8'd0;img500=8'd0;img501=8'd0;img502=8'd0;img503=8'd0;img504=8'd0;img505=8'd0;img506=8'd0;img507=8'd0;img508=8'd0;img509=8'd0;img510=8'd0;img511=8'd0;img512=8'd0;img513=8'd0;img514=8'd27;img515=8'd43;img516=8'd41;img517=8'd0;img518=8'd0;img519=8'd0;img520=8'd11;img521=8'd111;img522=8'd118;img523=8'd14;img524=8'd0;img525=8'd0;img526=8'd0;img527=8'd0;img528=8'd0;img529=8'd0;img530=8'd0;img531=8'd0;img532=8'd0;img533=8'd0;img534=8'd0;img535=8'd0;img536=8'd0;img537=8'd0;img538=8'd0;img539=8'd0;img540=8'd0;img541=8'd0;img542=8'd0;img543=8'd0;img544=8'd0;img545=8'd0;img546=8'd0;img547=8'd0;img548=8'd12;img549=8'd112;img550=8'd113;img551=8'd0;img552=8'd0;img553=8'd0;img554=8'd0;img555=8'd0;img556=8'd0;img557=8'd0;img558=8'd0;img559=8'd0;img560=8'd0;img561=8'd0;img562=8'd0;img563=8'd0;img564=8'd0;img565=8'd0;img566=8'd0;img567=8'd0;img568=8'd0;img569=8'd0;img570=8'd0;img571=8'd0;img572=8'd0;img573=8'd0;img574=8'd0;img575=8'd0;img576=8'd36;img577=8'd127;img578=8'd62;img579=8'd0;img580=8'd0;img581=8'd0;img582=8'd0;img583=8'd0;img584=8'd0;img585=8'd0;img586=8'd0;img587=8'd0;img588=8'd0;img589=8'd0;img590=8'd0;img591=8'd0;img592=8'd0;img593=8'd0;img594=8'd0;img595=8'd0;img596=8'd0;img597=8'd0;img598=8'd0;img599=8'd0;img600=8'd0;img601=8'd0;img602=8'd0;img603=8'd0;img604=8'd84;img605=8'd127;img606=8'd96;img607=8'd0;img608=8'd0;img609=8'd0;img610=8'd0;img611=8'd0;img612=8'd0;img613=8'd0;img614=8'd0;img615=8'd0;img616=8'd0;img617=8'd0;img618=8'd0;img619=8'd0;img620=8'd0;img621=8'd0;img622=8'd0;img623=8'd0;img624=8'd0;img625=8'd0;img626=8'd0;img627=8'd0;img628=8'd0;img629=8'd0;img630=8'd0;img631=8'd0;img632=8'd84;img633=8'd127;img634=8'd119;img635=8'd17;img636=8'd0;img637=8'd0;img638=8'd0;img639=8'd0;img640=8'd0;img641=8'd0;img642=8'd0;img643=8'd0;img644=8'd0;img645=8'd0;img646=8'd0;img647=8'd0;img648=8'd0;img649=8'd0;img650=8'd0;img651=8'd0;img652=8'd0;img653=8'd0;img654=8'd0;img655=8'd0;img656=8'd0;img657=8'd0;img658=8'd0;img659=8'd0;img660=8'd84;img661=8'd127;img662=8'd127;img663=8'd41;img664=8'd0;img665=8'd0;img666=8'd0;img667=8'd0;img668=8'd0;img669=8'd0;img670=8'd0;img671=8'd0;img672=8'd0;img673=8'd0;img674=8'd0;img675=8'd0;img676=8'd0;img677=8'd0;img678=8'd0;img679=8'd0;img680=8'd0;img681=8'd0;img682=8'd0;img683=8'd0;img684=8'd0;img685=8'd0;img686=8'd0;img687=8'd0;img688=8'd84;img689=8'd127;img690=8'd127;img691=8'd41;img692=8'd0;img693=8'd0;img694=8'd0;img695=8'd0;img696=8'd0;img697=8'd0;img698=8'd0;img699=8'd0;img700=8'd0;img701=8'd0;img702=8'd0;img703=8'd0;img704=8'd0;img705=8'd0;img706=8'd0;img707=8'd0;img708=8'd0;img709=8'd0;img710=8'd0;img711=8'd0;img712=8'd0;img713=8'd0;img714=8'd0;img715=8'd0;img716=8'd49;img717=8'd117;img718=8'd121;img719=8'd23;img720=8'd0;img721=8'd0;img722=8'd0;img723=8'd0;img724=8'd0;img725=8'd0;img726=8'd0;img727=8'd0;img728=8'd0;img729=8'd0;img730=8'd0;img731=8'd0;img732=8'd0;img733=8'd0;img734=8'd0;img735=8'd0;img736=8'd0;img737=8'd0;img738=8'd0;img739=8'd0;img740=8'd0;img741=8'd0;img742=8'd0;img743=8'd0;img744=8'd0;img745=8'd0;img746=8'd0;img747=8'd0;img748=8'd0;img749=8'd0;img750=8'd0;img751=8'd0;img752=8'd0;img753=8'd0;img754=8'd0;img755=8'd0;img756=8'd0;img757=8'd0;img758=8'd0;img759=8'd0;img760=8'd0;img761=8'd0;img762=8'd0;img763=8'd0;img764=8'd0;img765=8'd0;img766=8'd0;img767=8'd0;img768=8'd0;img769=8'd0;img770=8'd0;img771=8'd0;img772=8'd0;img773=8'd0;img774=8'd0;img775=8'd0;img776=8'd0;img777=8'd0;img778=8'd0;img779=8'd0;img780=8'd0;img781=8'd0;img782=8'd0;img783=8'd0;
$display("hit: %d :",hit);
#100 $finish;
end

endmodule 
