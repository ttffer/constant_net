`timescale 1ns / 1ps
module net
#(
DATAWIDTH=64,
BUFFCNT=2,
IMG_SZ=784
)
(
input clk,
input rst,
input  [7:0] img0,img1,img2,img3,img4,img5,img6,img7,img8,img9,img10,img11,img12,img13,img14,img15,img16,img17,img18,img19,img20,img21,img22,img23,img24,img25,img26,img27,img28,img29,img30,img31,img32,img33,img34,img35,img36,img37,img38,img39,img40,img41,img42,img43,img44,img45,img46,img47,img48,img49,img50,img51,img52,img53,img54,img55,img56,img57,img58,img59,img60,img61,img62,img63,img64,img65,img66,img67,img68,img69,img70,img71,img72,img73,img74,img75,img76,img77,img78,img79,img80,img81,img82,img83,img84,img85,img86,img87,img88,img89,img90,img91,img92,img93,img94,img95,img96,img97,img98,img99,img100,img101,img102,img103,img104,img105,img106,img107,img108,img109,img110,img111,img112,img113,img114,img115,img116,img117,img118,img119,img120,img121,img122,img123,img124,img125,img126,img127,img128,img129,img130,img131,img132,img133,img134,img135,img136,img137,img138,img139,img140,img141,img142,img143,img144,img145,img146,img147,img148,img149,img150,img151,img152,img153,img154,img155,img156,img157,img158,img159,img160,img161,img162,img163,img164,img165,img166,img167,img168,img169,img170,img171,img172,img173,img174,img175,img176,img177,img178,img179,img180,img181,img182,img183,img184,img185,img186,img187,img188,img189,img190,img191,img192,img193,img194,img195,img196,img197,img198,img199,img200,img201,img202,img203,img204,img205,img206,img207,img208,img209,img210,img211,img212,img213,img214,img215,img216,img217,img218,img219,img220,img221,img222,img223,img224,img225,img226,img227,img228,img229,img230,img231,img232,img233,img234,img235,img236,img237,img238,img239,img240,img241,img242,img243,img244,img245,img246,img247,img248,img249,img250,img251,img252,img253,img254,img255,img256,img257,img258,img259,img260,img261,img262,img263,img264,img265,img266,img267,img268,img269,img270,img271,img272,img273,img274,img275,img276,img277,img278,img279,img280,img281,img282,img283,img284,img285,img286,img287,img288,img289,img290,img291,img292,img293,img294,img295,img296,img297,img298,img299,img300,img301,img302,img303,img304,img305,img306,img307,img308,img309,img310,img311,img312,img313,img314,img315,img316,img317,img318,img319,img320,img321,img322,img323,img324,img325,img326,img327,img328,img329,img330,img331,img332,img333,img334,img335,img336,img337,img338,img339,img340,img341,img342,img343,img344,img345,img346,img347,img348,img349,img350,img351,img352,img353,img354,img355,img356,img357,img358,img359,img360,img361,img362,img363,img364,img365,img366,img367,img368,img369,img370,img371,img372,img373,img374,img375,img376,img377,img378,img379,img380,img381,img382,img383,img384,img385,img386,img387,img388,img389,img390,img391,img392,img393,img394,img395,img396,img397,img398,img399,img400,img401,img402,img403,img404,img405,img406,img407,img408,img409,img410,img411,img412,img413,img414,img415,img416,img417,img418,img419,img420,img421,img422,img423,img424,img425,img426,img427,img428,img429,img430,img431,img432,img433,img434,img435,img436,img437,img438,img439,img440,img441,img442,img443,img444,img445,img446,img447,img448,img449,img450,img451,img452,img453,img454,img455,img456,img457,img458,img459,img460,img461,img462,img463,img464,img465,img466,img467,img468,img469,img470,img471,img472,img473,img474,img475,img476,img477,img478,img479,img480,img481,img482,img483,img484,img485,img486,img487,img488,img489,img490,img491,img492,img493,img494,img495,img496,img497,img498,img499,img500,img501,img502,img503,img504,img505,img506,img507,img508,img509,img510,img511,img512,img513,img514,img515,img516,img517,img518,img519,img520,img521,img522,img523,img524,img525,img526,img527,img528,img529,img530,img531,img532,img533,img534,img535,img536,img537,img538,img539,img540,img541,img542,img543,img544,img545,img546,img547,img548,img549,img550,img551,img552,img553,img554,img555,img556,img557,img558,img559,img560,img561,img562,img563,img564,img565,img566,img567,img568,img569,img570,img571,img572,img573,img574,img575,img576,img577,img578,img579,img580,img581,img582,img583,img584,img585,img586,img587,img588,img589,img590,img591,img592,img593,img594,img595,img596,img597,img598,img599,img600,img601,img602,img603,img604,img605,img606,img607,img608,img609,img610,img611,img612,img613,img614,img615,img616,img617,img618,img619,img620,img621,img622,img623,img624,img625,img626,img627,img628,img629,img630,img631,img632,img633,img634,img635,img636,img637,img638,img639,img640,img641,img642,img643,img644,img645,img646,img647,img648,img649,img650,img651,img652,img653,img654,img655,img656,img657,img658,img659,img660,img661,img662,img663,img664,img665,img666,img667,img668,img669,img670,img671,img672,img673,img674,img675,img676,img677,img678,img679,img680,img681,img682,img683,img684,img685,img686,img687,img688,img689,img690,img691,img692,img693,img694,img695,img696,img697,img698,img699,img700,img701,img702,img703,img704,img705,img706,img707,img708,img709,img710,img711,img712,img713,img714,img715,img716,img717,img718,img719,img720,img721,img722,img723,img724,img725,img726,img727,img728,img729,img730,img731,img732,img733,img734,img735,img736,img737,img738,img739,img740,img741,img742,img743,img744,img745,img746,img747,img748,img749,img750,img751,img752,img753,img754,img755,img756,img757,img758,img759,img760,img761,img762,img763,img764,img765,img766,img767,img768,img769,img770,img771,img772,img773,img774,img775,img776,img777,img778,img779,img780,img781,img782,img783,

output    reg [4-1:0]predict

);
reg    [DATAWIDTH-1:0] in_buf  [0:783];
reg    [DATAWIDTH-1:0] result[0:9];
/////Start Declatation////////

wire [DATAWIDTH-1:0]   in_buf_weight00;
wire [DATAWIDTH-1:0]   in_buf_weight01;
wire [DATAWIDTH-1:0]   in_buf_weight02;
wire [DATAWIDTH-1:0]   in_buf_weight03;
wire [DATAWIDTH-1:0]   in_buf_weight04;
wire [DATAWIDTH-1:0]   in_buf_weight05;
wire [DATAWIDTH-1:0]   in_buf_weight06;
wire [DATAWIDTH-1:0]   in_buf_weight07;
wire [DATAWIDTH-1:0]   in_buf_weight08;
wire [DATAWIDTH-1:0]   in_buf_weight09;
wire [DATAWIDTH-1:0]   in_buf_weight010;
wire [DATAWIDTH-1:0]   in_buf_weight011;
wire [DATAWIDTH-1:0]   in_buf_weight012;
wire [DATAWIDTH-1:0]   in_buf_weight013;
wire [DATAWIDTH-1:0]   in_buf_weight014;
wire [DATAWIDTH-1:0]   in_buf_weight015;
wire [DATAWIDTH-1:0]   in_buf_weight016;
wire [DATAWIDTH-1:0]   in_buf_weight017;
wire [DATAWIDTH-1:0]   in_buf_weight018;
wire [DATAWIDTH-1:0]   in_buf_weight019;
wire [DATAWIDTH-1:0]   in_buf_weight020;
wire [DATAWIDTH-1:0]   in_buf_weight021;
wire [DATAWIDTH-1:0]   in_buf_weight022;
wire [DATAWIDTH-1:0]   in_buf_weight023;
wire [DATAWIDTH-1:0]   in_buf_weight024;
wire [DATAWIDTH-1:0]   in_buf_weight025;
wire [DATAWIDTH-1:0]   in_buf_weight026;
wire [DATAWIDTH-1:0]   in_buf_weight027;
wire [DATAWIDTH-1:0]   in_buf_weight028;
wire [DATAWIDTH-1:0]   in_buf_weight029;
wire [DATAWIDTH-1:0]   in_buf_weight030;
wire [DATAWIDTH-1:0]   in_buf_weight031;
wire [DATAWIDTH-1:0]   in_buf_weight032;
wire [DATAWIDTH-1:0]   in_buf_weight033;
wire [DATAWIDTH-1:0]   in_buf_weight034;
wire [DATAWIDTH-1:0]   in_buf_weight035;
wire [DATAWIDTH-1:0]   in_buf_weight036;
wire [DATAWIDTH-1:0]   in_buf_weight037;
wire [DATAWIDTH-1:0]   in_buf_weight038;
wire [DATAWIDTH-1:0]   in_buf_weight039;
wire [DATAWIDTH-1:0]   in_buf_weight040;
wire [DATAWIDTH-1:0]   in_buf_weight041;
wire [DATAWIDTH-1:0]   in_buf_weight042;
wire [DATAWIDTH-1:0]   in_buf_weight043;
wire [DATAWIDTH-1:0]   in_buf_weight044;
wire [DATAWIDTH-1:0]   in_buf_weight045;
wire [DATAWIDTH-1:0]   in_buf_weight046;
wire [DATAWIDTH-1:0]   in_buf_weight047;
wire [DATAWIDTH-1:0]   in_buf_weight048;
wire [DATAWIDTH-1:0]   in_buf_weight049;
wire [DATAWIDTH-1:0]   in_buf_weight050;
wire [DATAWIDTH-1:0]   in_buf_weight051;
wire [DATAWIDTH-1:0]   in_buf_weight052;
wire [DATAWIDTH-1:0]   in_buf_weight053;
wire [DATAWIDTH-1:0]   in_buf_weight054;
wire [DATAWIDTH-1:0]   in_buf_weight055;
wire [DATAWIDTH-1:0]   in_buf_weight056;
wire [DATAWIDTH-1:0]   in_buf_weight057;
wire [DATAWIDTH-1:0]   in_buf_weight058;
wire [DATAWIDTH-1:0]   in_buf_weight059;
wire [DATAWIDTH-1:0]   in_buf_weight060;
wire [DATAWIDTH-1:0]   in_buf_weight061;
wire [DATAWIDTH-1:0]   in_buf_weight062;
wire [DATAWIDTH-1:0]   in_buf_weight063;
assign in_buf_weight00=in_buf[0]*(-3)+in_buf[1]*(-2)+in_buf[2]*(-1)+in_buf[3]*(0)+in_buf[4]*(3)+in_buf[5]*(-3)+in_buf[6]*(0)+in_buf[7]*(0)+in_buf[8]*(0)+in_buf[9]*(1)+in_buf[10]*(-2)+in_buf[11]*(0)+in_buf[12]*(0)+in_buf[13]*(1)+in_buf[14]*(-9)+in_buf[15]*(-6)+in_buf[16]*(1)+in_buf[17]*(3)+in_buf[18]*(2)+in_buf[19]*(0)+in_buf[20]*(-2)+in_buf[21]*(-1)+in_buf[22]*(2)+in_buf[23]*(3)+in_buf[24]*(0)+in_buf[25]*(0)+in_buf[26]*(-1)+in_buf[27]*(3)+in_buf[28]*(1)+in_buf[29]*(-3)+in_buf[30]*(1)+in_buf[31]*(1)+in_buf[32]*(7)+in_buf[33]*(0)+in_buf[34]*(0)+in_buf[35]*(7)+in_buf[36]*(5)+in_buf[37]*(11)+in_buf[38]*(8)+in_buf[39]*(7)+in_buf[40]*(31)+in_buf[41]*(39)+in_buf[42]*(36)+in_buf[43]*(41)+in_buf[44]*(31)+in_buf[45]*(18)+in_buf[46]*(35)+in_buf[47]*(35)+in_buf[48]*(28)+in_buf[49]*(8)+in_buf[50]*(3)+in_buf[51]*(1)+in_buf[52]*(0)+in_buf[53]*(4)+in_buf[54]*(-1)+in_buf[55]*(0)+in_buf[56]*(-3)+in_buf[57]*(0)+in_buf[58]*(22)+in_buf[59]*(7)+in_buf[60]*(20)+in_buf[61]*(1)+in_buf[62]*(0)+in_buf[63]*(9)+in_buf[64]*(-10)+in_buf[65]*(-29)+in_buf[66]*(-35)+in_buf[67]*(-5)+in_buf[68]*(-12)+in_buf[69]*(10)+in_buf[70]*(6)+in_buf[71]*(14)+in_buf[72]*(2)+in_buf[73]*(7)+in_buf[74]*(21)+in_buf[75]*(25)+in_buf[76]*(21)+in_buf[77]*(18)+in_buf[78]*(32)+in_buf[79]*(34)+in_buf[80]*(-12)+in_buf[81]*(-4)+in_buf[82]*(0)+in_buf[83]*(0)+in_buf[84]*(-1)+in_buf[85]*(2)+in_buf[86]*(30)+in_buf[87]*(21)+in_buf[88]*(22)+in_buf[89]*(-17)+in_buf[90]*(-14)+in_buf[91]*(0)+in_buf[92]*(-34)+in_buf[93]*(-28)+in_buf[94]*(-49)+in_buf[95]*(-44)+in_buf[96]*(-14)+in_buf[97]*(3)+in_buf[98]*(14)+in_buf[99]*(3)+in_buf[100]*(-10)+in_buf[101]*(13)+in_buf[102]*(17)+in_buf[103]*(31)+in_buf[104]*(32)+in_buf[105]*(19)+in_buf[106]*(21)+in_buf[107]*(1)+in_buf[108]*(2)+in_buf[109]*(-7)+in_buf[110]*(17)+in_buf[111]*(0)+in_buf[112]*(-3)+in_buf[113]*(-8)+in_buf[114]*(16)+in_buf[115]*(-3)+in_buf[116]*(-28)+in_buf[117]*(-27)+in_buf[118]*(-48)+in_buf[119]*(-60)+in_buf[120]*(-64)+in_buf[121]*(-46)+in_buf[122]*(-14)+in_buf[123]*(-17)+in_buf[124]*(-5)+in_buf[125]*(12)+in_buf[126]*(-7)+in_buf[127]*(0)+in_buf[128]*(0)+in_buf[129]*(-1)+in_buf[130]*(1)+in_buf[131]*(3)+in_buf[132]*(-2)+in_buf[133]*(5)+in_buf[134]*(-1)+in_buf[135]*(6)+in_buf[136]*(-25)+in_buf[137]*(3)+in_buf[138]*(0)+in_buf[139]*(5)+in_buf[140]*(3)+in_buf[141]*(4)+in_buf[142]*(36)+in_buf[143]*(-4)+in_buf[144]*(-26)+in_buf[145]*(-40)+in_buf[146]*(-72)+in_buf[147]*(-65)+in_buf[148]*(-39)+in_buf[149]*(-20)+in_buf[150]*(0)+in_buf[151]*(5)+in_buf[152]*(4)+in_buf[153]*(9)+in_buf[154]*(10)+in_buf[155]*(2)+in_buf[156]*(-2)+in_buf[157]*(-7)+in_buf[158]*(2)+in_buf[159]*(-5)+in_buf[160]*(1)+in_buf[161]*(2)+in_buf[162]*(-5)+in_buf[163]*(6)+in_buf[164]*(-5)+in_buf[165]*(21)+in_buf[166]*(5)+in_buf[167]*(-4)+in_buf[168]*(3)+in_buf[169]*(-19)+in_buf[170]*(15)+in_buf[171]*(-12)+in_buf[172]*(-34)+in_buf[173]*(-38)+in_buf[174]*(-70)+in_buf[175]*(-44)+in_buf[176]*(-22)+in_buf[177]*(-17)+in_buf[178]*(0)+in_buf[179]*(14)+in_buf[180]*(6)+in_buf[181]*(12)+in_buf[182]*(6)+in_buf[183]*(-2)+in_buf[184]*(-16)+in_buf[185]*(-14)+in_buf[186]*(2)+in_buf[187]*(6)+in_buf[188]*(14)+in_buf[189]*(-5)+in_buf[190]*(2)+in_buf[191]*(-9)+in_buf[192]*(29)+in_buf[193]*(51)+in_buf[194]*(4)+in_buf[195]*(3)+in_buf[196]*(4)+in_buf[197]*(-28)+in_buf[198]*(-5)+in_buf[199]*(-38)+in_buf[200]*(-70)+in_buf[201]*(-51)+in_buf[202]*(-47)+in_buf[203]*(-23)+in_buf[204]*(-6)+in_buf[205]*(8)+in_buf[206]*(4)+in_buf[207]*(8)+in_buf[208]*(16)+in_buf[209]*(11)+in_buf[210]*(14)+in_buf[211]*(4)+in_buf[212]*(6)+in_buf[213]*(10)+in_buf[214]*(19)+in_buf[215]*(14)+in_buf[216]*(30)+in_buf[217]*(19)+in_buf[218]*(16)+in_buf[219]*(9)+in_buf[220]*(4)+in_buf[221]*(10)+in_buf[222]*(29)+in_buf[223]*(22)+in_buf[224]*(-2)+in_buf[225]*(-26)+in_buf[226]*(-22)+in_buf[227]*(-47)+in_buf[228]*(-62)+in_buf[229]*(-45)+in_buf[230]*(-15)+in_buf[231]*(-16)+in_buf[232]*(-18)+in_buf[233]*(-1)+in_buf[234]*(-3)+in_buf[235]*(12)+in_buf[236]*(16)+in_buf[237]*(16)+in_buf[238]*(24)+in_buf[239]*(13)+in_buf[240]*(7)+in_buf[241]*(13)+in_buf[242]*(15)+in_buf[243]*(20)+in_buf[244]*(36)+in_buf[245]*(25)+in_buf[246]*(19)+in_buf[247]*(23)+in_buf[248]*(33)+in_buf[249]*(30)+in_buf[250]*(33)+in_buf[251]*(27)+in_buf[252]*(3)+in_buf[253]*(-1)+in_buf[254]*(-34)+in_buf[255]*(-42)+in_buf[256]*(-25)+in_buf[257]*(-21)+in_buf[258]*(-12)+in_buf[259]*(-15)+in_buf[260]*(-12)+in_buf[261]*(-18)+in_buf[262]*(-3)+in_buf[263]*(12)+in_buf[264]*(7)+in_buf[265]*(27)+in_buf[266]*(32)+in_buf[267]*(3)+in_buf[268]*(-16)+in_buf[269]*(-11)+in_buf[270]*(7)+in_buf[271]*(9)+in_buf[272]*(4)+in_buf[273]*(16)+in_buf[274]*(12)+in_buf[275]*(9)+in_buf[276]*(32)+in_buf[277]*(31)+in_buf[278]*(24)+in_buf[279]*(25)+in_buf[280]*(4)+in_buf[281]*(7)+in_buf[282]*(-21)+in_buf[283]*(-38)+in_buf[284]*(-12)+in_buf[285]*(-19)+in_buf[286]*(-18)+in_buf[287]*(-1)+in_buf[288]*(-6)+in_buf[289]*(-1)+in_buf[290]*(6)+in_buf[291]*(8)+in_buf[292]*(14)+in_buf[293]*(30)+in_buf[294]*(1)+in_buf[295]*(-34)+in_buf[296]*(-57)+in_buf[297]*(-53)+in_buf[298]*(-45)+in_buf[299]*(-36)+in_buf[300]*(-29)+in_buf[301]*(-30)+in_buf[302]*(-31)+in_buf[303]*(-46)+in_buf[304]*(-22)+in_buf[305]*(34)+in_buf[306]*(47)+in_buf[307]*(4)+in_buf[308]*(2)+in_buf[309]*(5)+in_buf[310]*(-3)+in_buf[311]*(-45)+in_buf[312]*(-18)+in_buf[313]*(-2)+in_buf[314]*(-7)+in_buf[315]*(-4)+in_buf[316]*(-13)+in_buf[317]*(-15)+in_buf[318]*(8)+in_buf[319]*(-4)+in_buf[320]*(3)+in_buf[321]*(-2)+in_buf[322]*(-34)+in_buf[323]*(-56)+in_buf[324]*(-44)+in_buf[325]*(-45)+in_buf[326]*(-59)+in_buf[327]*(-82)+in_buf[328]*(-99)+in_buf[329]*(-82)+in_buf[330]*(-77)+in_buf[331]*(-83)+in_buf[332]*(-65)+in_buf[333]*(14)+in_buf[334]*(33)+in_buf[335]*(29)+in_buf[336]*(9)+in_buf[337]*(-2)+in_buf[338]*(7)+in_buf[339]*(-21)+in_buf[340]*(-26)+in_buf[341]*(-7)+in_buf[342]*(0)+in_buf[343]*(-3)+in_buf[344]*(-3)+in_buf[345]*(-11)+in_buf[346]*(14)+in_buf[347]*(6)+in_buf[348]*(12)+in_buf[349]*(6)+in_buf[350]*(-14)+in_buf[351]*(-24)+in_buf[352]*(-18)+in_buf[353]*(-30)+in_buf[354]*(-23)+in_buf[355]*(-75)+in_buf[356]*(-92)+in_buf[357]*(-102)+in_buf[358]*(-99)+in_buf[359]*(-106)+in_buf[360]*(-81)+in_buf[361]*(-31)+in_buf[362]*(0)+in_buf[363]*(38)+in_buf[364]*(0)+in_buf[365]*(2)+in_buf[366]*(8)+in_buf[367]*(-18)+in_buf[368]*(-7)+in_buf[369]*(9)+in_buf[370]*(17)+in_buf[371]*(12)+in_buf[372]*(-12)+in_buf[373]*(-2)+in_buf[374]*(5)+in_buf[375]*(8)+in_buf[376]*(16)+in_buf[377]*(5)+in_buf[378]*(2)+in_buf[379]*(7)+in_buf[380]*(0)+in_buf[381]*(-2)+in_buf[382]*(3)+in_buf[383]*(6)+in_buf[384]*(-22)+in_buf[385]*(-42)+in_buf[386]*(-73)+in_buf[387]*(-76)+in_buf[388]*(-73)+in_buf[389]*(-33)+in_buf[390]*(-8)+in_buf[391]*(-2)+in_buf[392]*(16)+in_buf[393]*(-14)+in_buf[394]*(-7)+in_buf[395]*(-20)+in_buf[396]*(6)+in_buf[397]*(9)+in_buf[398]*(25)+in_buf[399]*(23)+in_buf[400]*(0)+in_buf[401]*(8)+in_buf[402]*(8)+in_buf[403]*(-1)+in_buf[404]*(-3)+in_buf[405]*(-8)+in_buf[406]*(-1)+in_buf[407]*(7)+in_buf[408]*(4)+in_buf[409]*(7)+in_buf[410]*(12)+in_buf[411]*(1)+in_buf[412]*(3)+in_buf[413]*(-17)+in_buf[414]*(-22)+in_buf[415]*(-4)+in_buf[416]*(-5)+in_buf[417]*(-13)+in_buf[418]*(-37)+in_buf[419]*(2)+in_buf[420]*(11)+in_buf[421]*(-11)+in_buf[422]*(-1)+in_buf[423]*(5)+in_buf[424]*(3)+in_buf[425]*(15)+in_buf[426]*(10)+in_buf[427]*(19)+in_buf[428]*(7)+in_buf[429]*(11)+in_buf[430]*(9)+in_buf[431]*(1)+in_buf[432]*(10)+in_buf[433]*(-6)+in_buf[434]*(-13)+in_buf[435]*(-5)+in_buf[436]*(9)+in_buf[437]*(17)+in_buf[438]*(16)+in_buf[439]*(-12)+in_buf[440]*(0)+in_buf[441]*(2)+in_buf[442]*(-24)+in_buf[443]*(10)+in_buf[444]*(11)+in_buf[445]*(22)+in_buf[446]*(-33)+in_buf[447]*(-23)+in_buf[448]*(-1)+in_buf[449]*(-10)+in_buf[450]*(-25)+in_buf[451]*(21)+in_buf[452]*(-7)+in_buf[453]*(5)+in_buf[454]*(-9)+in_buf[455]*(5)+in_buf[456]*(9)+in_buf[457]*(0)+in_buf[458]*(1)+in_buf[459]*(6)+in_buf[460]*(0)+in_buf[461]*(-7)+in_buf[462]*(5)+in_buf[463]*(11)+in_buf[464]*(2)+in_buf[465]*(25)+in_buf[466]*(14)+in_buf[467]*(4)+in_buf[468]*(9)+in_buf[469]*(1)+in_buf[470]*(0)+in_buf[471]*(-14)+in_buf[472]*(11)+in_buf[473]*(26)+in_buf[474]*(-26)+in_buf[475]*(-25)+in_buf[476]*(0)+in_buf[477]*(-8)+in_buf[478]*(-1)+in_buf[479]*(13)+in_buf[480]*(-1)+in_buf[481]*(11)+in_buf[482]*(16)+in_buf[483]*(20)+in_buf[484]*(0)+in_buf[485]*(-9)+in_buf[486]*(-1)+in_buf[487]*(-7)+in_buf[488]*(-3)+in_buf[489]*(-6)+in_buf[490]*(8)+in_buf[491]*(22)+in_buf[492]*(3)+in_buf[493]*(19)+in_buf[494]*(28)+in_buf[495]*(8)+in_buf[496]*(10)+in_buf[497]*(1)+in_buf[498]*(5)+in_buf[499]*(6)+in_buf[500]*(1)+in_buf[501]*(-9)+in_buf[502]*(-26)+in_buf[503]*(-29)+in_buf[504]*(-2)+in_buf[505]*(-5)+in_buf[506]*(-6)+in_buf[507]*(-3)+in_buf[508]*(5)+in_buf[509]*(8)+in_buf[510]*(23)+in_buf[511]*(21)+in_buf[512]*(4)+in_buf[513]*(-6)+in_buf[514]*(-34)+in_buf[515]*(-19)+in_buf[516]*(0)+in_buf[517]*(-7)+in_buf[518]*(10)+in_buf[519]*(23)+in_buf[520]*(9)+in_buf[521]*(8)+in_buf[522]*(9)+in_buf[523]*(3)+in_buf[524]*(12)+in_buf[525]*(3)+in_buf[526]*(-16)+in_buf[527]*(3)+in_buf[528]*(7)+in_buf[529]*(4)+in_buf[530]*(-38)+in_buf[531]*(-42)+in_buf[532]*(3)+in_buf[533]*(-8)+in_buf[534]*(17)+in_buf[535]*(-16)+in_buf[536]*(2)+in_buf[537]*(0)+in_buf[538]*(31)+in_buf[539]*(10)+in_buf[540]*(7)+in_buf[541]*(6)+in_buf[542]*(-22)+in_buf[543]*(-7)+in_buf[544]*(5)+in_buf[545]*(-6)+in_buf[546]*(17)+in_buf[547]*(21)+in_buf[548]*(9)+in_buf[549]*(-1)+in_buf[550]*(10)+in_buf[551]*(9)+in_buf[552]*(10)+in_buf[553]*(-6)+in_buf[554]*(-12)+in_buf[555]*(16)+in_buf[556]*(33)+in_buf[557]*(11)+in_buf[558]*(-40)+in_buf[559]*(-28)+in_buf[560]*(3)+in_buf[561]*(-14)+in_buf[562]*(17)+in_buf[563]*(-25)+in_buf[564]*(-4)+in_buf[565]*(2)+in_buf[566]*(10)+in_buf[567]*(-6)+in_buf[568]*(11)+in_buf[569]*(14)+in_buf[570]*(-4)+in_buf[571]*(-5)+in_buf[572]*(2)+in_buf[573]*(-4)+in_buf[574]*(4)+in_buf[575]*(12)+in_buf[576]*(9)+in_buf[577]*(11)+in_buf[578]*(16)+in_buf[579]*(20)+in_buf[580]*(3)+in_buf[581]*(-6)+in_buf[582]*(5)+in_buf[583]*(14)+in_buf[584]*(19)+in_buf[585]*(15)+in_buf[586]*(-32)+in_buf[587]*(3)+in_buf[588]*(4)+in_buf[589]*(-16)+in_buf[590]*(-31)+in_buf[591]*(-29)+in_buf[592]*(19)+in_buf[593]*(13)+in_buf[594]*(4)+in_buf[595]*(-6)+in_buf[596]*(0)+in_buf[597]*(13)+in_buf[598]*(8)+in_buf[599]*(6)+in_buf[600]*(2)+in_buf[601]*(0)+in_buf[602]*(20)+in_buf[603]*(16)+in_buf[604]*(7)+in_buf[605]*(4)+in_buf[606]*(20)+in_buf[607]*(15)+in_buf[608]*(25)+in_buf[609]*(12)+in_buf[610]*(4)+in_buf[611]*(3)+in_buf[612]*(6)+in_buf[613]*(27)+in_buf[614]*(20)+in_buf[615]*(-4)+in_buf[616]*(2)+in_buf[617]*(-21)+in_buf[618]*(-46)+in_buf[619]*(18)+in_buf[620]*(10)+in_buf[621]*(11)+in_buf[622]*(-13)+in_buf[623]*(-14)+in_buf[624]*(-11)+in_buf[625]*(-2)+in_buf[626]*(3)+in_buf[627]*(5)+in_buf[628]*(7)+in_buf[629]*(-4)+in_buf[630]*(4)+in_buf[631]*(20)+in_buf[632]*(12)+in_buf[633]*(8)+in_buf[634]*(9)+in_buf[635]*(4)+in_buf[636]*(15)+in_buf[637]*(7)+in_buf[638]*(-18)+in_buf[639]*(14)+in_buf[640]*(1)+in_buf[641]*(12)+in_buf[642]*(28)+in_buf[643]*(0)+in_buf[644]*(2)+in_buf[645]*(0)+in_buf[646]*(-27)+in_buf[647]*(22)+in_buf[648]*(28)+in_buf[649]*(20)+in_buf[650]*(16)+in_buf[651]*(-14)+in_buf[652]*(-10)+in_buf[653]*(2)+in_buf[654]*(5)+in_buf[655]*(1)+in_buf[656]*(7)+in_buf[657]*(-4)+in_buf[658]*(10)+in_buf[659]*(13)+in_buf[660]*(-5)+in_buf[661]*(-1)+in_buf[662]*(-11)+in_buf[663]*(0)+in_buf[664]*(2)+in_buf[665]*(-5)+in_buf[666]*(-3)+in_buf[667]*(9)+in_buf[668]*(9)+in_buf[669]*(17)+in_buf[670]*(31)+in_buf[671]*(2)+in_buf[672]*(2)+in_buf[673]*(-1)+in_buf[674]*(-34)+in_buf[675]*(-1)+in_buf[676]*(-16)+in_buf[677]*(-10)+in_buf[678]*(16)+in_buf[679]*(20)+in_buf[680]*(-3)+in_buf[681]*(8)+in_buf[682]*(4)+in_buf[683]*(-3)+in_buf[684]*(0)+in_buf[685]*(7)+in_buf[686]*(4)+in_buf[687]*(2)+in_buf[688]*(2)+in_buf[689]*(21)+in_buf[690]*(26)+in_buf[691]*(-7)+in_buf[692]*(-9)+in_buf[693]*(-9)+in_buf[694]*(2)+in_buf[695]*(-13)+in_buf[696]*(10)+in_buf[697]*(15)+in_buf[698]*(24)+in_buf[699]*(4)+in_buf[700]*(0)+in_buf[701]*(-1)+in_buf[702]*(1)+in_buf[703]*(6)+in_buf[704]*(-4)+in_buf[705]*(-22)+in_buf[706]*(-1)+in_buf[707]*(17)+in_buf[708]*(2)+in_buf[709]*(24)+in_buf[710]*(1)+in_buf[711]*(7)+in_buf[712]*(18)+in_buf[713]*(0)+in_buf[714]*(-9)+in_buf[715]*(1)+in_buf[716]*(-2)+in_buf[717]*(7)+in_buf[718]*(11)+in_buf[719]*(30)+in_buf[720]*(37)+in_buf[721]*(37)+in_buf[722]*(48)+in_buf[723]*(37)+in_buf[724]*(25)+in_buf[725]*(2)+in_buf[726]*(5)+in_buf[727]*(-3)+in_buf[728]*(0)+in_buf[729]*(2)+in_buf[730]*(3)+in_buf[731]*(-2)+in_buf[732]*(1)+in_buf[733]*(-1)+in_buf[734]*(-18)+in_buf[735]*(-13)+in_buf[736]*(-8)+in_buf[737]*(26)+in_buf[738]*(9)+in_buf[739]*(-28)+in_buf[740]*(-18)+in_buf[741]*(-6)+in_buf[742]*(-13)+in_buf[743]*(9)+in_buf[744]*(15)+in_buf[745]*(-20)+in_buf[746]*(-8)+in_buf[747]*(10)+in_buf[748]*(9)+in_buf[749]*(22)+in_buf[750]*(25)+in_buf[751]*(4)+in_buf[752]*(3)+in_buf[753]*(0)+in_buf[754]*(0)+in_buf[755]*(3)+in_buf[756]*(1)+in_buf[757]*(-3)+in_buf[758]*(-1)+in_buf[759]*(2)+in_buf[760]*(-1)+in_buf[761]*(2)+in_buf[762]*(-3)+in_buf[763]*(-8)+in_buf[764]*(-11)+in_buf[765]*(-11)+in_buf[766]*(-9)+in_buf[767]*(3)+in_buf[768]*(-2)+in_buf[769]*(5)+in_buf[770]*(-12)+in_buf[771]*(6)+in_buf[772]*(-3)+in_buf[773]*(-23)+in_buf[774]*(-25)+in_buf[775]*(-20)+in_buf[776]*(-6)+in_buf[777]*(-7)+in_buf[778]*(0)+in_buf[779]*(3)+in_buf[780]*(4)+in_buf[781]*(-3)+in_buf[782]*(2)+in_buf[783]*(2);
assign in_buf_weight01=in_buf[0]*(-3)+in_buf[1]*(0)+in_buf[2]*(-2)+in_buf[3]*(-3)+in_buf[4]*(0)+in_buf[5]*(3)+in_buf[6]*(-3)+in_buf[7]*(1)+in_buf[8]*(4)+in_buf[9]*(3)+in_buf[10]*(3)+in_buf[11]*(4)+in_buf[12]*(10)+in_buf[13]*(3)+in_buf[14]*(-21)+in_buf[15]*(-17)+in_buf[16]*(-2)+in_buf[17]*(3)+in_buf[18]*(1)+in_buf[19]*(-2)+in_buf[20]*(-2)+in_buf[21]*(-2)+in_buf[22]*(0)+in_buf[23]*(-3)+in_buf[24]*(-3)+in_buf[25]*(2)+in_buf[26]*(4)+in_buf[27]*(-3)+in_buf[28]*(1)+in_buf[29]*(4)+in_buf[30]*(0)+in_buf[31]*(3)+in_buf[32]*(-5)+in_buf[33]*(4)+in_buf[34]*(8)+in_buf[35]*(9)+in_buf[36]*(11)+in_buf[37]*(6)+in_buf[38]*(23)+in_buf[39]*(0)+in_buf[40]*(-9)+in_buf[41]*(-18)+in_buf[42]*(14)+in_buf[43]*(-16)+in_buf[44]*(-28)+in_buf[45]*(-22)+in_buf[46]*(31)+in_buf[47]*(28)+in_buf[48]*(25)+in_buf[49]*(9)+in_buf[50]*(0)+in_buf[51]*(0)+in_buf[52]*(-3)+in_buf[53]*(-2)+in_buf[54]*(0)+in_buf[55]*(0)+in_buf[56]*(3)+in_buf[57]*(-1)+in_buf[58]*(0)+in_buf[59]*(-8)+in_buf[60]*(-8)+in_buf[61]*(13)+in_buf[62]*(24)+in_buf[63]*(19)+in_buf[64]*(3)+in_buf[65]*(6)+in_buf[66]*(31)+in_buf[67]*(28)+in_buf[68]*(51)+in_buf[69]*(69)+in_buf[70]*(53)+in_buf[71]*(55)+in_buf[72]*(15)+in_buf[73]*(15)+in_buf[74]*(-2)+in_buf[75]*(25)+in_buf[76]*(19)+in_buf[77]*(14)+in_buf[78]*(30)+in_buf[79]*(12)+in_buf[80]*(34)+in_buf[81]*(-3)+in_buf[82]*(4)+in_buf[83]*(0)+in_buf[84]*(-1)+in_buf[85]*(1)+in_buf[86]*(7)+in_buf[87]*(-9)+in_buf[88]*(-8)+in_buf[89]*(1)+in_buf[90]*(23)+in_buf[91]*(11)+in_buf[92]*(-8)+in_buf[93]*(8)+in_buf[94]*(-3)+in_buf[95]*(17)+in_buf[96]*(14)+in_buf[97]*(28)+in_buf[98]*(-6)+in_buf[99]*(4)+in_buf[100]*(18)+in_buf[101]*(0)+in_buf[102]*(-9)+in_buf[103]*(-9)+in_buf[104]*(-24)+in_buf[105]*(8)+in_buf[106]*(21)+in_buf[107]*(25)+in_buf[108]*(-11)+in_buf[109]*(-24)+in_buf[110]*(-9)+in_buf[111]*(-1)+in_buf[112]*(3)+in_buf[113]*(1)+in_buf[114]*(8)+in_buf[115]*(-26)+in_buf[116]*(11)+in_buf[117]*(46)+in_buf[118]*(47)+in_buf[119]*(33)+in_buf[120]*(44)+in_buf[121]*(30)+in_buf[122]*(27)+in_buf[123]*(11)+in_buf[124]*(14)+in_buf[125]*(24)+in_buf[126]*(8)+in_buf[127]*(2)+in_buf[128]*(11)+in_buf[129]*(-6)+in_buf[130]*(-23)+in_buf[131]*(-10)+in_buf[132]*(-4)+in_buf[133]*(0)+in_buf[134]*(18)+in_buf[135]*(6)+in_buf[136]*(0)+in_buf[137]*(-30)+in_buf[138]*(-34)+in_buf[139]*(-1)+in_buf[140]*(1)+in_buf[141]*(0)+in_buf[142]*(10)+in_buf[143]*(26)+in_buf[144]*(48)+in_buf[145]*(43)+in_buf[146]*(36)+in_buf[147]*(24)+in_buf[148]*(1)+in_buf[149]*(-11)+in_buf[150]*(-7)+in_buf[151]*(-16)+in_buf[152]*(3)+in_buf[153]*(-2)+in_buf[154]*(4)+in_buf[155]*(14)+in_buf[156]*(-1)+in_buf[157]*(-13)+in_buf[158]*(-8)+in_buf[159]*(-2)+in_buf[160]*(7)+in_buf[161]*(7)+in_buf[162]*(16)+in_buf[163]*(12)+in_buf[164]*(15)+in_buf[165]*(0)+in_buf[166]*(-34)+in_buf[167]*(15)+in_buf[168]*(-1)+in_buf[169]*(-10)+in_buf[170]*(-27)+in_buf[171]*(20)+in_buf[172]*(6)+in_buf[173]*(-17)+in_buf[174]*(-6)+in_buf[175]*(-12)+in_buf[176]*(-26)+in_buf[177]*(-25)+in_buf[178]*(-2)+in_buf[179]*(-1)+in_buf[180]*(-16)+in_buf[181]*(-12)+in_buf[182]*(-15)+in_buf[183]*(0)+in_buf[184]*(-1)+in_buf[185]*(-15)+in_buf[186]*(-2)+in_buf[187]*(-8)+in_buf[188]*(9)+in_buf[189]*(11)+in_buf[190]*(1)+in_buf[191]*(13)+in_buf[192]*(-8)+in_buf[193]*(5)+in_buf[194]*(-17)+in_buf[195]*(14)+in_buf[196]*(2)+in_buf[197]*(-22)+in_buf[198]*(-37)+in_buf[199]*(-9)+in_buf[200]*(18)+in_buf[201]*(-8)+in_buf[202]*(-13)+in_buf[203]*(-23)+in_buf[204]*(-49)+in_buf[205]*(-27)+in_buf[206]*(-18)+in_buf[207]*(-9)+in_buf[208]*(-2)+in_buf[209]*(1)+in_buf[210]*(-1)+in_buf[211]*(-1)+in_buf[212]*(-5)+in_buf[213]*(0)+in_buf[214]*(-2)+in_buf[215]*(-3)+in_buf[216]*(5)+in_buf[217]*(11)+in_buf[218]*(18)+in_buf[219]*(13)+in_buf[220]*(7)+in_buf[221]*(-9)+in_buf[222]*(-2)+in_buf[223]*(-7)+in_buf[224]*(-33)+in_buf[225]*(-29)+in_buf[226]*(4)+in_buf[227]*(8)+in_buf[228]*(17)+in_buf[229]*(4)+in_buf[230]*(-25)+in_buf[231]*(-31)+in_buf[232]*(-46)+in_buf[233]*(-38)+in_buf[234]*(-11)+in_buf[235]*(-7)+in_buf[236]*(-2)+in_buf[237]*(10)+in_buf[238]*(-2)+in_buf[239]*(4)+in_buf[240]*(-3)+in_buf[241]*(9)+in_buf[242]*(0)+in_buf[243]*(2)+in_buf[244]*(-2)+in_buf[245]*(8)+in_buf[246]*(0)+in_buf[247]*(0)+in_buf[248]*(2)+in_buf[249]*(-6)+in_buf[250]*(19)+in_buf[251]*(-14)+in_buf[252]*(-20)+in_buf[253]*(-37)+in_buf[254]*(26)+in_buf[255]*(20)+in_buf[256]*(8)+in_buf[257]*(-8)+in_buf[258]*(-30)+in_buf[259]*(-32)+in_buf[260]*(-32)+in_buf[261]*(-11)+in_buf[262]*(1)+in_buf[263]*(4)+in_buf[264]*(9)+in_buf[265]*(15)+in_buf[266]*(4)+in_buf[267]*(3)+in_buf[268]*(1)+in_buf[269]*(0)+in_buf[270]*(0)+in_buf[271]*(-4)+in_buf[272]*(2)+in_buf[273]*(15)+in_buf[274]*(-5)+in_buf[275]*(-16)+in_buf[276]*(0)+in_buf[277]*(-23)+in_buf[278]*(10)+in_buf[279]*(-11)+in_buf[280]*(-22)+in_buf[281]*(-15)+in_buf[282]*(-15)+in_buf[283]*(8)+in_buf[284]*(5)+in_buf[285]*(-10)+in_buf[286]*(-37)+in_buf[287]*(-38)+in_buf[288]*(-29)+in_buf[289]*(-24)+in_buf[290]*(2)+in_buf[291]*(9)+in_buf[292]*(20)+in_buf[293]*(-3)+in_buf[294]*(-3)+in_buf[295]*(-7)+in_buf[296]*(-7)+in_buf[297]*(0)+in_buf[298]*(-2)+in_buf[299]*(-5)+in_buf[300]*(-15)+in_buf[301]*(1)+in_buf[302]*(-21)+in_buf[303]*(-21)+in_buf[304]*(-31)+in_buf[305]*(-19)+in_buf[306]*(-10)+in_buf[307]*(-11)+in_buf[308]*(-20)+in_buf[309]*(-36)+in_buf[310]*(-23)+in_buf[311]*(-4)+in_buf[312]*(21)+in_buf[313]*(6)+in_buf[314]*(-20)+in_buf[315]*(-8)+in_buf[316]*(-15)+in_buf[317]*(3)+in_buf[318]*(13)+in_buf[319]*(12)+in_buf[320]*(6)+in_buf[321]*(-12)+in_buf[322]*(-9)+in_buf[323]*(0)+in_buf[324]*(5)+in_buf[325]*(0)+in_buf[326]*(1)+in_buf[327]*(0)+in_buf[328]*(-3)+in_buf[329]*(-2)+in_buf[330]*(-20)+in_buf[331]*(-26)+in_buf[332]*(-22)+in_buf[333]*(-21)+in_buf[334]*(-15)+in_buf[335]*(-28)+in_buf[336]*(-3)+in_buf[337]*(-12)+in_buf[338]*(-18)+in_buf[339]*(-2)+in_buf[340]*(25)+in_buf[341]*(9)+in_buf[342]*(5)+in_buf[343]*(9)+in_buf[344]*(11)+in_buf[345]*(22)+in_buf[346]*(10)+in_buf[347]*(5)+in_buf[348]*(0)+in_buf[349]*(-12)+in_buf[350]*(0)+in_buf[351]*(-1)+in_buf[352]*(16)+in_buf[353]*(22)+in_buf[354]*(12)+in_buf[355]*(5)+in_buf[356]*(-13)+in_buf[357]*(-5)+in_buf[358]*(-4)+in_buf[359]*(-17)+in_buf[360]*(-33)+in_buf[361]*(-31)+in_buf[362]*(-40)+in_buf[363]*(-35)+in_buf[364]*(22)+in_buf[365]*(4)+in_buf[366]*(-22)+in_buf[367]*(-16)+in_buf[368]*(21)+in_buf[369]*(6)+in_buf[370]*(15)+in_buf[371]*(15)+in_buf[372]*(26)+in_buf[373]*(20)+in_buf[374]*(11)+in_buf[375]*(0)+in_buf[376]*(-11)+in_buf[377]*(-3)+in_buf[378]*(5)+in_buf[379]*(13)+in_buf[380]*(19)+in_buf[381]*(33)+in_buf[382]*(21)+in_buf[383]*(-1)+in_buf[384]*(-15)+in_buf[385]*(0)+in_buf[386]*(-2)+in_buf[387]*(-11)+in_buf[388]*(-33)+in_buf[389]*(-19)+in_buf[390]*(-29)+in_buf[391]*(-7)+in_buf[392]*(-17)+in_buf[393]*(7)+in_buf[394]*(11)+in_buf[395]*(5)+in_buf[396]*(21)+in_buf[397]*(21)+in_buf[398]*(12)+in_buf[399]*(24)+in_buf[400]*(24)+in_buf[401]*(17)+in_buf[402]*(-2)+in_buf[403]*(-15)+in_buf[404]*(-14)+in_buf[405]*(1)+in_buf[406]*(12)+in_buf[407]*(16)+in_buf[408]*(36)+in_buf[409]*(18)+in_buf[410]*(7)+in_buf[411]*(-6)+in_buf[412]*(-16)+in_buf[413]*(-2)+in_buf[414]*(1)+in_buf[415]*(-26)+in_buf[416]*(-48)+in_buf[417]*(2)+in_buf[418]*(1)+in_buf[419]*(-6)+in_buf[420]*(-17)+in_buf[421]*(0)+in_buf[422]*(48)+in_buf[423]*(25)+in_buf[424]*(24)+in_buf[425]*(8)+in_buf[426]*(-10)+in_buf[427]*(12)+in_buf[428]*(27)+in_buf[429]*(22)+in_buf[430]*(10)+in_buf[431]*(-8)+in_buf[432]*(-11)+in_buf[433]*(20)+in_buf[434]*(21)+in_buf[435]*(24)+in_buf[436]*(32)+in_buf[437]*(-4)+in_buf[438]*(-16)+in_buf[439]*(-9)+in_buf[440]*(-30)+in_buf[441]*(-28)+in_buf[442]*(7)+in_buf[443]*(-28)+in_buf[444]*(-50)+in_buf[445]*(11)+in_buf[446]*(34)+in_buf[447]*(15)+in_buf[448]*(0)+in_buf[449]*(10)+in_buf[450]*(32)+in_buf[451]*(-2)+in_buf[452]*(15)+in_buf[453]*(0)+in_buf[454]*(8)+in_buf[455]*(29)+in_buf[456]*(18)+in_buf[457]*(11)+in_buf[458]*(12)+in_buf[459]*(-7)+in_buf[460]*(-6)+in_buf[461]*(4)+in_buf[462]*(18)+in_buf[463]*(19)+in_buf[464]*(15)+in_buf[465]*(-13)+in_buf[466]*(-16)+in_buf[467]*(-18)+in_buf[468]*(-28)+in_buf[469]*(-8)+in_buf[470]*(0)+in_buf[471]*(-2)+in_buf[472]*(-9)+in_buf[473]*(24)+in_buf[474]*(4)+in_buf[475]*(14)+in_buf[476]*(0)+in_buf[477]*(1)+in_buf[478]*(41)+in_buf[479]*(0)+in_buf[480]*(12)+in_buf[481]*(-4)+in_buf[482]*(-11)+in_buf[483]*(14)+in_buf[484]*(18)+in_buf[485]*(0)+in_buf[486]*(0)+in_buf[487]*(-12)+in_buf[488]*(-3)+in_buf[489]*(0)+in_buf[490]*(22)+in_buf[491]*(17)+in_buf[492]*(-10)+in_buf[493]*(-28)+in_buf[494]*(-20)+in_buf[495]*(-13)+in_buf[496]*(-16)+in_buf[497]*(15)+in_buf[498]*(10)+in_buf[499]*(8)+in_buf[500]*(12)+in_buf[501]*(35)+in_buf[502]*(41)+in_buf[503]*(10)+in_buf[504]*(-27)+in_buf[505]*(2)+in_buf[506]*(25)+in_buf[507]*(23)+in_buf[508]*(12)+in_buf[509]*(-4)+in_buf[510]*(-9)+in_buf[511]*(10)+in_buf[512]*(9)+in_buf[513]*(4)+in_buf[514]*(-19)+in_buf[515]*(-20)+in_buf[516]*(-22)+in_buf[517]*(-7)+in_buf[518]*(16)+in_buf[519]*(6)+in_buf[520]*(-10)+in_buf[521]*(-15)+in_buf[522]*(-4)+in_buf[523]*(-1)+in_buf[524]*(4)+in_buf[525]*(22)+in_buf[526]*(41)+in_buf[527]*(37)+in_buf[528]*(23)+in_buf[529]*(44)+in_buf[530]*(36)+in_buf[531]*(31)+in_buf[532]*(10)+in_buf[533]*(-38)+in_buf[534]*(-7)+in_buf[535]*(16)+in_buf[536]*(12)+in_buf[537]*(-7)+in_buf[538]*(-11)+in_buf[539]*(9)+in_buf[540]*(0)+in_buf[541]*(-8)+in_buf[542]*(-18)+in_buf[543]*(-23)+in_buf[544]*(-38)+in_buf[545]*(-19)+in_buf[546]*(2)+in_buf[547]*(25)+in_buf[548]*(29)+in_buf[549]*(3)+in_buf[550]*(6)+in_buf[551]*(10)+in_buf[552]*(4)+in_buf[553]*(39)+in_buf[554]*(37)+in_buf[555]*(30)+in_buf[556]*(22)+in_buf[557]*(26)+in_buf[558]*(45)+in_buf[559]*(9)+in_buf[560]*(0)+in_buf[561]*(-8)+in_buf[562]*(-4)+in_buf[563]*(16)+in_buf[564]*(14)+in_buf[565]*(-11)+in_buf[566]*(6)+in_buf[567]*(10)+in_buf[568]*(-8)+in_buf[569]*(-5)+in_buf[570]*(-11)+in_buf[571]*(-12)+in_buf[572]*(-14)+in_buf[573]*(-15)+in_buf[574]*(10)+in_buf[575]*(21)+in_buf[576]*(36)+in_buf[577]*(23)+in_buf[578]*(41)+in_buf[579]*(32)+in_buf[580]*(30)+in_buf[581]*(38)+in_buf[582]*(31)+in_buf[583]*(32)+in_buf[584]*(25)+in_buf[585]*(11)+in_buf[586]*(43)+in_buf[587]*(2)+in_buf[588]*(3)+in_buf[589]*(8)+in_buf[590]*(-2)+in_buf[591]*(16)+in_buf[592]*(-4)+in_buf[593]*(0)+in_buf[594]*(17)+in_buf[595]*(10)+in_buf[596]*(14)+in_buf[597]*(0)+in_buf[598]*(3)+in_buf[599]*(-16)+in_buf[600]*(-12)+in_buf[601]*(1)+in_buf[602]*(5)+in_buf[603]*(12)+in_buf[604]*(14)+in_buf[605]*(14)+in_buf[606]*(33)+in_buf[607]*(31)+in_buf[608]*(31)+in_buf[609]*(15)+in_buf[610]*(16)+in_buf[611]*(17)+in_buf[612]*(9)+in_buf[613]*(-3)+in_buf[614]*(-25)+in_buf[615]*(3)+in_buf[616]*(8)+in_buf[617]*(10)+in_buf[618]*(7)+in_buf[619]*(7)+in_buf[620]*(-3)+in_buf[621]*(18)+in_buf[622]*(12)+in_buf[623]*(6)+in_buf[624]*(7)+in_buf[625]*(0)+in_buf[626]*(-4)+in_buf[627]*(-10)+in_buf[628]*(-13)+in_buf[629]*(-7)+in_buf[630]*(-13)+in_buf[631]*(-1)+in_buf[632]*(-17)+in_buf[633]*(-4)+in_buf[634]*(28)+in_buf[635]*(29)+in_buf[636]*(18)+in_buf[637]*(22)+in_buf[638]*(9)+in_buf[639]*(-2)+in_buf[640]*(3)+in_buf[641]*(-12)+in_buf[642]*(-15)+in_buf[643]*(-5)+in_buf[644]*(4)+in_buf[645]*(-2)+in_buf[646]*(-9)+in_buf[647]*(0)+in_buf[648]*(-33)+in_buf[649]*(-14)+in_buf[650]*(4)+in_buf[651]*(-5)+in_buf[652]*(-4)+in_buf[653]*(-10)+in_buf[654]*(-19)+in_buf[655]*(-31)+in_buf[656]*(-16)+in_buf[657]*(-15)+in_buf[658]*(-10)+in_buf[659]*(-3)+in_buf[660]*(-11)+in_buf[661]*(-4)+in_buf[662]*(20)+in_buf[663]*(13)+in_buf[664]*(17)+in_buf[665]*(13)+in_buf[666]*(10)+in_buf[667]*(-2)+in_buf[668]*(-8)+in_buf[669]*(-13)+in_buf[670]*(0)+in_buf[671]*(0)+in_buf[672]*(-1)+in_buf[673]*(2)+in_buf[674]*(-1)+in_buf[675]*(-30)+in_buf[676]*(-21)+in_buf[677]*(-28)+in_buf[678]*(-5)+in_buf[679]*(3)+in_buf[680]*(8)+in_buf[681]*(17)+in_buf[682]*(-11)+in_buf[683]*(-20)+in_buf[684]*(-18)+in_buf[685]*(-13)+in_buf[686]*(-9)+in_buf[687]*(-20)+in_buf[688]*(-29)+in_buf[689]*(-10)+in_buf[690]*(4)+in_buf[691]*(2)+in_buf[692]*(-8)+in_buf[693]*(22)+in_buf[694]*(22)+in_buf[695]*(1)+in_buf[696]*(2)+in_buf[697]*(22)+in_buf[698]*(26)+in_buf[699]*(3)+in_buf[700]*(-1)+in_buf[701]*(-1)+in_buf[702]*(34)+in_buf[703]*(-34)+in_buf[704]*(-39)+in_buf[705]*(-42)+in_buf[706]*(-8)+in_buf[707]*(-1)+in_buf[708]*(30)+in_buf[709]*(16)+in_buf[710]*(-9)+in_buf[711]*(4)+in_buf[712]*(20)+in_buf[713]*(-12)+in_buf[714]*(3)+in_buf[715]*(-9)+in_buf[716]*(-33)+in_buf[717]*(-32)+in_buf[718]*(-6)+in_buf[719]*(-18)+in_buf[720]*(-3)+in_buf[721]*(16)+in_buf[722]*(2)+in_buf[723]*(-11)+in_buf[724]*(-27)+in_buf[725]*(17)+in_buf[726]*(19)+in_buf[727]*(1)+in_buf[728]*(4)+in_buf[729]*(3)+in_buf[730]*(3)+in_buf[731]*(13)+in_buf[732]*(25)+in_buf[733]*(1)+in_buf[734]*(6)+in_buf[735]*(-2)+in_buf[736]*(-2)+in_buf[737]*(-17)+in_buf[738]*(15)+in_buf[739]*(16)+in_buf[740]*(7)+in_buf[741]*(-18)+in_buf[742]*(5)+in_buf[743]*(21)+in_buf[744]*(9)+in_buf[745]*(-13)+in_buf[746]*(-12)+in_buf[747]*(-39)+in_buf[748]*(-14)+in_buf[749]*(9)+in_buf[750]*(0)+in_buf[751]*(16)+in_buf[752]*(20)+in_buf[753]*(-7)+in_buf[754]*(4)+in_buf[755]*(3)+in_buf[756]*(-1)+in_buf[757]*(3)+in_buf[758]*(4)+in_buf[759]*(0)+in_buf[760]*(-19)+in_buf[761]*(-29)+in_buf[762]*(6)+in_buf[763]*(15)+in_buf[764]*(7)+in_buf[765]*(6)+in_buf[766]*(5)+in_buf[767]*(15)+in_buf[768]*(15)+in_buf[769]*(4)+in_buf[770]*(5)+in_buf[771]*(23)+in_buf[772]*(-4)+in_buf[773]*(-13)+in_buf[774]*(5)+in_buf[775]*(27)+in_buf[776]*(37)+in_buf[777]*(4)+in_buf[778]*(5)+in_buf[779]*(-16)+in_buf[780]*(4)+in_buf[781]*(4)+in_buf[782]*(0)+in_buf[783]*(0);
assign in_buf_weight02=in_buf[0]*(4)+in_buf[1]*(-1)+in_buf[2]*(4)+in_buf[3]*(1)+in_buf[4]*(-1)+in_buf[5]*(2)+in_buf[6]*(4)+in_buf[7]*(0)+in_buf[8]*(3)+in_buf[9]*(-3)+in_buf[10]*(3)+in_buf[11]*(0)+in_buf[12]*(10)+in_buf[13]*(15)+in_buf[14]*(19)+in_buf[15]*(11)+in_buf[16]*(-3)+in_buf[17]*(-2)+in_buf[18]*(-1)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(2)+in_buf[22]*(0)+in_buf[23]*(0)+in_buf[24]*(-1)+in_buf[25]*(2)+in_buf[26]*(-3)+in_buf[27]*(0)+in_buf[28]*(2)+in_buf[29]*(4)+in_buf[30]*(-1)+in_buf[31]*(-1)+in_buf[32]*(4)+in_buf[33]*(8)+in_buf[34]*(11)+in_buf[35]*(11)+in_buf[36]*(15)+in_buf[37]*(15)+in_buf[38]*(30)+in_buf[39]*(10)+in_buf[40]*(11)+in_buf[41]*(4)+in_buf[42]*(-19)+in_buf[43]*(-7)+in_buf[44]*(-10)+in_buf[45]*(15)+in_buf[46]*(33)+in_buf[47]*(31)+in_buf[48]*(32)+in_buf[49]*(25)+in_buf[50]*(20)+in_buf[51]*(13)+in_buf[52]*(0)+in_buf[53]*(0)+in_buf[54]*(0)+in_buf[55]*(0)+in_buf[56]*(-1)+in_buf[57]*(-3)+in_buf[58]*(21)+in_buf[59]*(3)+in_buf[60]*(16)+in_buf[61]*(10)+in_buf[62]*(15)+in_buf[63]*(22)+in_buf[64]*(40)+in_buf[65]*(31)+in_buf[66]*(17)+in_buf[67]*(41)+in_buf[68]*(28)+in_buf[69]*(-2)+in_buf[70]*(22)+in_buf[71]*(4)+in_buf[72]*(-2)+in_buf[73]*(27)+in_buf[74]*(20)+in_buf[75]*(8)+in_buf[76]*(-5)+in_buf[77]*(0)+in_buf[78]*(9)+in_buf[79]*(2)+in_buf[80]*(0)+in_buf[81]*(-2)+in_buf[82]*(0)+in_buf[83]*(-2)+in_buf[84]*(-1)+in_buf[85]*(3)+in_buf[86]*(-13)+in_buf[87]*(-3)+in_buf[88]*(8)+in_buf[89]*(21)+in_buf[90]*(32)+in_buf[91]*(-1)+in_buf[92]*(-2)+in_buf[93]*(24)+in_buf[94]*(0)+in_buf[95]*(11)+in_buf[96]*(8)+in_buf[97]*(-1)+in_buf[98]*(1)+in_buf[99]*(-6)+in_buf[100]*(10)+in_buf[101]*(9)+in_buf[102]*(-2)+in_buf[103]*(7)+in_buf[104]*(3)+in_buf[105]*(11)+in_buf[106]*(5)+in_buf[107]*(-9)+in_buf[108]*(3)+in_buf[109]*(-6)+in_buf[110]*(6)+in_buf[111]*(-3)+in_buf[112]*(3)+in_buf[113]*(0)+in_buf[114]*(-18)+in_buf[115]*(-17)+in_buf[116]*(35)+in_buf[117]*(27)+in_buf[118]*(24)+in_buf[119]*(-6)+in_buf[120]*(6)+in_buf[121]*(6)+in_buf[122]*(2)+in_buf[123]*(6)+in_buf[124]*(10)+in_buf[125]*(-1)+in_buf[126]*(3)+in_buf[127]*(-20)+in_buf[128]*(0)+in_buf[129]*(12)+in_buf[130]*(-11)+in_buf[131]*(-2)+in_buf[132]*(-8)+in_buf[133]*(-23)+in_buf[134]*(-37)+in_buf[135]*(-38)+in_buf[136]*(-28)+in_buf[137]*(-35)+in_buf[138]*(-7)+in_buf[139]*(3)+in_buf[140]*(0)+in_buf[141]*(0)+in_buf[142]*(8)+in_buf[143]*(-8)+in_buf[144]*(24)+in_buf[145]*(8)+in_buf[146]*(11)+in_buf[147]*(3)+in_buf[148]*(24)+in_buf[149]*(21)+in_buf[150]*(25)+in_buf[151]*(9)+in_buf[152]*(10)+in_buf[153]*(-10)+in_buf[154]*(-5)+in_buf[155]*(-9)+in_buf[156]*(4)+in_buf[157]*(-25)+in_buf[158]*(-34)+in_buf[159]*(-20)+in_buf[160]*(-6)+in_buf[161]*(-16)+in_buf[162]*(-45)+in_buf[163]*(-29)+in_buf[164]*(-23)+in_buf[165]*(-31)+in_buf[166]*(-16)+in_buf[167]*(1)+in_buf[168]*(2)+in_buf[169]*(-1)+in_buf[170]*(3)+in_buf[171]*(6)+in_buf[172]*(28)+in_buf[173]*(22)+in_buf[174]*(0)+in_buf[175]*(3)+in_buf[176]*(21)+in_buf[177]*(29)+in_buf[178]*(21)+in_buf[179]*(36)+in_buf[180]*(15)+in_buf[181]*(-4)+in_buf[182]*(-13)+in_buf[183]*(-15)+in_buf[184]*(-25)+in_buf[185]*(-22)+in_buf[186]*(-49)+in_buf[187]*(-35)+in_buf[188]*(-25)+in_buf[189]*(-21)+in_buf[190]*(-16)+in_buf[191]*(-9)+in_buf[192]*(8)+in_buf[193]*(-5)+in_buf[194]*(-22)+in_buf[195]*(10)+in_buf[196]*(6)+in_buf[197]*(4)+in_buf[198]*(30)+in_buf[199]*(2)+in_buf[200]*(2)+in_buf[201]*(6)+in_buf[202]*(1)+in_buf[203]*(0)+in_buf[204]*(23)+in_buf[205]*(30)+in_buf[206]*(42)+in_buf[207]*(26)+in_buf[208]*(6)+in_buf[209]*(-12)+in_buf[210]*(-30)+in_buf[211]*(-24)+in_buf[212]*(-26)+in_buf[213]*(-17)+in_buf[214]*(-20)+in_buf[215]*(-30)+in_buf[216]*(-20)+in_buf[217]*(-3)+in_buf[218]*(-19)+in_buf[219]*(-24)+in_buf[220]*(5)+in_buf[221]*(9)+in_buf[222]*(-7)+in_buf[223]*(-2)+in_buf[224]*(12)+in_buf[225]*(-8)+in_buf[226]*(31)+in_buf[227]*(-25)+in_buf[228]*(6)+in_buf[229]*(-5)+in_buf[230]*(4)+in_buf[231]*(4)+in_buf[232]*(16)+in_buf[233]*(38)+in_buf[234]*(36)+in_buf[235]*(14)+in_buf[236]*(7)+in_buf[237]*(-17)+in_buf[238]*(-14)+in_buf[239]*(-12)+in_buf[240]*(-23)+in_buf[241]*(-22)+in_buf[242]*(-22)+in_buf[243]*(-15)+in_buf[244]*(-2)+in_buf[245]*(-2)+in_buf[246]*(-10)+in_buf[247]*(8)+in_buf[248]*(-12)+in_buf[249]*(-4)+in_buf[250]*(13)+in_buf[251]*(-29)+in_buf[252]*(8)+in_buf[253]*(15)+in_buf[254]*(-11)+in_buf[255]*(-44)+in_buf[256]*(-1)+in_buf[257]*(-6)+in_buf[258]*(-26)+in_buf[259]*(-12)+in_buf[260]*(4)+in_buf[261]*(13)+in_buf[262]*(4)+in_buf[263]*(8)+in_buf[264]*(7)+in_buf[265]*(-8)+in_buf[266]*(-18)+in_buf[267]*(-20)+in_buf[268]*(-17)+in_buf[269]*(-10)+in_buf[270]*(-5)+in_buf[271]*(-2)+in_buf[272]*(6)+in_buf[273]*(7)+in_buf[274]*(8)+in_buf[275]*(10)+in_buf[276]*(1)+in_buf[277]*(-15)+in_buf[278]*(-5)+in_buf[279]*(18)+in_buf[280]*(8)+in_buf[281]*(5)+in_buf[282]*(-22)+in_buf[283]*(-32)+in_buf[284]*(-10)+in_buf[285]*(-8)+in_buf[286]*(-17)+in_buf[287]*(-11)+in_buf[288]*(1)+in_buf[289]*(1)+in_buf[290]*(-2)+in_buf[291]*(-5)+in_buf[292]*(-7)+in_buf[293]*(-4)+in_buf[294]*(-23)+in_buf[295]*(-20)+in_buf[296]*(1)+in_buf[297]*(10)+in_buf[298]*(0)+in_buf[299]*(-4)+in_buf[300]*(-4)+in_buf[301]*(3)+in_buf[302]*(3)+in_buf[303]*(1)+in_buf[304]*(21)+in_buf[305]*(-18)+in_buf[306]*(-25)+in_buf[307]*(0)+in_buf[308]*(5)+in_buf[309]*(36)+in_buf[310]*(-25)+in_buf[311]*(-5)+in_buf[312]*(-25)+in_buf[313]*(-23)+in_buf[314]*(-20)+in_buf[315]*(-18)+in_buf[316]*(-1)+in_buf[317]*(-1)+in_buf[318]*(-10)+in_buf[319]*(-2)+in_buf[320]*(5)+in_buf[321]*(-21)+in_buf[322]*(-26)+in_buf[323]*(-13)+in_buf[324]*(0)+in_buf[325]*(5)+in_buf[326]*(0)+in_buf[327]*(2)+in_buf[328]*(7)+in_buf[329]*(17)+in_buf[330]*(18)+in_buf[331]*(10)+in_buf[332]*(7)+in_buf[333]*(0)+in_buf[334]*(-32)+in_buf[335]*(-24)+in_buf[336]*(-2)+in_buf[337]*(-1)+in_buf[338]*(-32)+in_buf[339]*(-41)+in_buf[340]*(-44)+in_buf[341]*(-35)+in_buf[342]*(-36)+in_buf[343]*(-17)+in_buf[344]*(-5)+in_buf[345]*(-14)+in_buf[346]*(-7)+in_buf[347]*(4)+in_buf[348]*(15)+in_buf[349]*(-5)+in_buf[350]*(-5)+in_buf[351]*(-2)+in_buf[352]*(8)+in_buf[353]*(7)+in_buf[354]*(8)+in_buf[355]*(17)+in_buf[356]*(4)+in_buf[357]*(19)+in_buf[358]*(23)+in_buf[359]*(2)+in_buf[360]*(29)+in_buf[361]*(-5)+in_buf[362]*(-35)+in_buf[363]*(-33)+in_buf[364]*(-17)+in_buf[365]*(-3)+in_buf[366]*(-3)+in_buf[367]*(-36)+in_buf[368]*(-58)+in_buf[369]*(-3)+in_buf[370]*(-11)+in_buf[371]*(-19)+in_buf[372]*(-14)+in_buf[373]*(-14)+in_buf[374]*(0)+in_buf[375]*(-2)+in_buf[376]*(8)+in_buf[377]*(9)+in_buf[378]*(-3)+in_buf[379]*(6)+in_buf[380]*(6)+in_buf[381]*(2)+in_buf[382]*(15)+in_buf[383]*(13)+in_buf[384]*(8)+in_buf[385]*(20)+in_buf[386]*(11)+in_buf[387]*(28)+in_buf[388]*(13)+in_buf[389]*(-5)+in_buf[390]*(-9)+in_buf[391]*(9)+in_buf[392]*(-4)+in_buf[393]*(-2)+in_buf[394]*(5)+in_buf[395]*(-16)+in_buf[396]*(-46)+in_buf[397]*(-6)+in_buf[398]*(6)+in_buf[399]*(-11)+in_buf[400]*(0)+in_buf[401]*(-3)+in_buf[402]*(-2)+in_buf[403]*(5)+in_buf[404]*(4)+in_buf[405]*(9)+in_buf[406]*(10)+in_buf[407]*(6)+in_buf[408]*(17)+in_buf[409]*(8)+in_buf[410]*(15)+in_buf[411]*(16)+in_buf[412]*(1)+in_buf[413]*(20)+in_buf[414]*(32)+in_buf[415]*(24)+in_buf[416]*(6)+in_buf[417]*(20)+in_buf[418]*(10)+in_buf[419]*(20)+in_buf[420]*(-2)+in_buf[421]*(-1)+in_buf[422]*(-22)+in_buf[423]*(-17)+in_buf[424]*(-31)+in_buf[425]*(-9)+in_buf[426]*(6)+in_buf[427]*(10)+in_buf[428]*(2)+in_buf[429]*(-1)+in_buf[430]*(-14)+in_buf[431]*(-2)+in_buf[432]*(8)+in_buf[433]*(14)+in_buf[434]*(23)+in_buf[435]*(16)+in_buf[436]*(12)+in_buf[437]*(11)+in_buf[438]*(15)+in_buf[439]*(17)+in_buf[440]*(6)+in_buf[441]*(12)+in_buf[442]*(17)+in_buf[443]*(13)+in_buf[444]*(16)+in_buf[445]*(46)+in_buf[446]*(-17)+in_buf[447]*(40)+in_buf[448]*(3)+in_buf[449]*(0)+in_buf[450]*(-8)+in_buf[451]*(-31)+in_buf[452]*(-35)+in_buf[453]*(-2)+in_buf[454]*(13)+in_buf[455]*(-3)+in_buf[456]*(7)+in_buf[457]*(-4)+in_buf[458]*(-3)+in_buf[459]*(0)+in_buf[460]*(-1)+in_buf[461]*(6)+in_buf[462]*(16)+in_buf[463]*(7)+in_buf[464]*(19)+in_buf[465]*(23)+in_buf[466]*(9)+in_buf[467]*(2)+in_buf[468]*(-11)+in_buf[469]*(8)+in_buf[470]*(8)+in_buf[471]*(19)+in_buf[472]*(35)+in_buf[473]*(45)+in_buf[474]*(16)+in_buf[475]*(28)+in_buf[476]*(-2)+in_buf[477]*(-5)+in_buf[478]*(-12)+in_buf[479]*(-26)+in_buf[480]*(-26)+in_buf[481]*(-17)+in_buf[482]*(-11)+in_buf[483]*(-17)+in_buf[484]*(0)+in_buf[485]*(-16)+in_buf[486]*(-14)+in_buf[487]*(-3)+in_buf[488]*(13)+in_buf[489]*(18)+in_buf[490]*(17)+in_buf[491]*(6)+in_buf[492]*(16)+in_buf[493]*(13)+in_buf[494]*(11)+in_buf[495]*(5)+in_buf[496]*(8)+in_buf[497]*(4)+in_buf[498]*(13)+in_buf[499]*(25)+in_buf[500]*(27)+in_buf[501]*(46)+in_buf[502]*(13)+in_buf[503]*(18)+in_buf[504]*(-33)+in_buf[505]*(-8)+in_buf[506]*(-18)+in_buf[507]*(22)+in_buf[508]*(-21)+in_buf[509]*(-14)+in_buf[510]*(-7)+in_buf[511]*(4)+in_buf[512]*(-8)+in_buf[513]*(-26)+in_buf[514]*(-30)+in_buf[515]*(-4)+in_buf[516]*(30)+in_buf[517]*(26)+in_buf[518]*(20)+in_buf[519]*(12)+in_buf[520]*(0)+in_buf[521]*(6)+in_buf[522]*(5)+in_buf[523]*(-3)+in_buf[524]*(-14)+in_buf[525]*(-9)+in_buf[526]*(3)+in_buf[527]*(29)+in_buf[528]*(28)+in_buf[529]*(54)+in_buf[530]*(34)+in_buf[531]*(32)+in_buf[532]*(-16)+in_buf[533]*(-29)+in_buf[534]*(-22)+in_buf[535]*(26)+in_buf[536]*(-4)+in_buf[537]*(-5)+in_buf[538]*(-19)+in_buf[539]*(-13)+in_buf[540]*(-26)+in_buf[541]*(-31)+in_buf[542]*(-6)+in_buf[543]*(33)+in_buf[544]*(24)+in_buf[545]*(18)+in_buf[546]*(25)+in_buf[547]*(8)+in_buf[548]*(-6)+in_buf[549]*(6)+in_buf[550]*(5)+in_buf[551]*(-11)+in_buf[552]*(-4)+in_buf[553]*(-14)+in_buf[554]*(7)+in_buf[555]*(22)+in_buf[556]*(0)+in_buf[557]*(17)+in_buf[558]*(56)+in_buf[559]*(12)+in_buf[560]*(1)+in_buf[561]*(0)+in_buf[562]*(-1)+in_buf[563]*(1)+in_buf[564]*(-20)+in_buf[565]*(23)+in_buf[566]*(-20)+in_buf[567]*(-12)+in_buf[568]*(-39)+in_buf[569]*(-25)+in_buf[570]*(8)+in_buf[571]*(35)+in_buf[572]*(41)+in_buf[573]*(26)+in_buf[574]*(21)+in_buf[575]*(17)+in_buf[576]*(-17)+in_buf[577]*(-9)+in_buf[578]*(-6)+in_buf[579]*(-11)+in_buf[580]*(-3)+in_buf[581]*(-14)+in_buf[582]*(-4)+in_buf[583]*(-15)+in_buf[584]*(-5)+in_buf[585]*(-2)+in_buf[586]*(45)+in_buf[587]*(-5)+in_buf[588]*(-7)+in_buf[589]*(0)+in_buf[590]*(-6)+in_buf[591]*(-3)+in_buf[592]*(-30)+in_buf[593]*(0)+in_buf[594]*(-14)+in_buf[595]*(-31)+in_buf[596]*(-14)+in_buf[597]*(0)+in_buf[598]*(16)+in_buf[599]*(19)+in_buf[600]*(21)+in_buf[601]*(23)+in_buf[602]*(19)+in_buf[603]*(-7)+in_buf[604]*(-8)+in_buf[605]*(-1)+in_buf[606]*(-1)+in_buf[607]*(-1)+in_buf[608]*(-13)+in_buf[609]*(-27)+in_buf[610]*(-10)+in_buf[611]*(-11)+in_buf[612]*(-20)+in_buf[613]*(-1)+in_buf[614]*(48)+in_buf[615]*(5)+in_buf[616]*(-4)+in_buf[617]*(-11)+in_buf[618]*(-6)+in_buf[619]*(-32)+in_buf[620]*(-30)+in_buf[621]*(-17)+in_buf[622]*(-21)+in_buf[623]*(-11)+in_buf[624]*(-8)+in_buf[625]*(3)+in_buf[626]*(6)+in_buf[627]*(6)+in_buf[628]*(7)+in_buf[629]*(9)+in_buf[630]*(-3)+in_buf[631]*(-4)+in_buf[632]*(-12)+in_buf[633]*(-30)+in_buf[634]*(-33)+in_buf[635]*(-9)+in_buf[636]*(-23)+in_buf[637]*(-19)+in_buf[638]*(-7)+in_buf[639]*(-23)+in_buf[640]*(-36)+in_buf[641]*(-10)+in_buf[642]*(-17)+in_buf[643]*(0)+in_buf[644]*(-2)+in_buf[645]*(-3)+in_buf[646]*(-4)+in_buf[647]*(-34)+in_buf[648]*(-40)+in_buf[649]*(-20)+in_buf[650]*(-6)+in_buf[651]*(1)+in_buf[652]*(-2)+in_buf[653]*(-5)+in_buf[654]*(-20)+in_buf[655]*(-11)+in_buf[656]*(10)+in_buf[657]*(-3)+in_buf[658]*(5)+in_buf[659]*(-4)+in_buf[660]*(-16)+in_buf[661]*(-33)+in_buf[662]*(-26)+in_buf[663]*(-23)+in_buf[664]*(-27)+in_buf[665]*(3)+in_buf[666]*(10)+in_buf[667]*(-14)+in_buf[668]*(-38)+in_buf[669]*(-1)+in_buf[670]*(-21)+in_buf[671]*(-1)+in_buf[672]*(-2)+in_buf[673]*(0)+in_buf[674]*(4)+in_buf[675]*(-10)+in_buf[676]*(-22)+in_buf[677]*(-22)+in_buf[678]*(-20)+in_buf[679]*(-38)+in_buf[680]*(-20)+in_buf[681]*(-8)+in_buf[682]*(-20)+in_buf[683]*(-7)+in_buf[684]*(13)+in_buf[685]*(14)+in_buf[686]*(31)+in_buf[687]*(9)+in_buf[688]*(6)+in_buf[689]*(-22)+in_buf[690]*(-31)+in_buf[691]*(-39)+in_buf[692]*(-31)+in_buf[693]*(14)+in_buf[694]*(30)+in_buf[695]*(-17)+in_buf[696]*(39)+in_buf[697]*(12)+in_buf[698]*(0)+in_buf[699]*(0)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(-26)+in_buf[703]*(0)+in_buf[704]*(-29)+in_buf[705]*(-25)+in_buf[706]*(-7)+in_buf[707]*(-11)+in_buf[708]*(-17)+in_buf[709]*(0)+in_buf[710]*(-1)+in_buf[711]*(10)+in_buf[712]*(4)+in_buf[713]*(2)+in_buf[714]*(8)+in_buf[715]*(17)+in_buf[716]*(26)+in_buf[717]*(5)+in_buf[718]*(-30)+in_buf[719]*(-52)+in_buf[720]*(-39)+in_buf[721]*(-17)+in_buf[722]*(-4)+in_buf[723]*(-26)+in_buf[724]*(-34)+in_buf[725]*(-11)+in_buf[726]*(-1)+in_buf[727]*(4)+in_buf[728]*(1)+in_buf[729]*(0)+in_buf[730]*(1)+in_buf[731]*(0)+in_buf[732]*(-36)+in_buf[733]*(-34)+in_buf[734]*(-41)+in_buf[735]*(-33)+in_buf[736]*(-4)+in_buf[737]*(4)+in_buf[738]*(-15)+in_buf[739]*(-18)+in_buf[740]*(-11)+in_buf[741]*(-16)+in_buf[742]*(-29)+in_buf[743]*(9)+in_buf[744]*(1)+in_buf[745]*(-20)+in_buf[746]*(-25)+in_buf[747]*(-24)+in_buf[748]*(-34)+in_buf[749]*(-30)+in_buf[750]*(-38)+in_buf[751]*(-22)+in_buf[752]*(7)+in_buf[753]*(20)+in_buf[754]*(0)+in_buf[755]*(0)+in_buf[756]*(-1)+in_buf[757]*(2)+in_buf[758]*(-2)+in_buf[759]*(0)+in_buf[760]*(24)+in_buf[761]*(18)+in_buf[762]*(18)+in_buf[763]*(10)+in_buf[764]*(10)+in_buf[765]*(23)+in_buf[766]*(-21)+in_buf[767]*(-7)+in_buf[768]*(-1)+in_buf[769]*(-5)+in_buf[770]*(-59)+in_buf[771]*(10)+in_buf[772]*(29)+in_buf[773]*(5)+in_buf[774]*(3)+in_buf[775]*(1)+in_buf[776]*(1)+in_buf[777]*(2)+in_buf[778]*(-2)+in_buf[779]*(5)+in_buf[780]*(1)+in_buf[781]*(-1)+in_buf[782]*(2)+in_buf[783]*(3);
assign in_buf_weight03=in_buf[0]*(0)+in_buf[1]*(-3)+in_buf[2]*(3)+in_buf[3]*(0)+in_buf[4]*(4)+in_buf[5]*(2)+in_buf[6]*(1)+in_buf[7]*(0)+in_buf[8]*(0)+in_buf[9]*(0)+in_buf[10]*(0)+in_buf[11]*(3)+in_buf[12]*(6)+in_buf[13]*(6)+in_buf[14]*(0)+in_buf[15]*(3)+in_buf[16]*(1)+in_buf[17]*(4)+in_buf[18]*(3)+in_buf[19]*(0)+in_buf[20]*(4)+in_buf[21]*(2)+in_buf[22]*(-2)+in_buf[23]*(-1)+in_buf[24]*(0)+in_buf[25]*(-3)+in_buf[26]*(3)+in_buf[27]*(1)+in_buf[28]*(2)+in_buf[29]*(-2)+in_buf[30]*(-2)+in_buf[31]*(2)+in_buf[32]*(9)+in_buf[33]*(6)+in_buf[34]*(13)+in_buf[35]*(15)+in_buf[36]*(12)+in_buf[37]*(12)+in_buf[38]*(6)+in_buf[39]*(0)+in_buf[40]*(9)+in_buf[41]*(8)+in_buf[42]*(-13)+in_buf[43]*(37)+in_buf[44]*(30)+in_buf[45]*(41)+in_buf[46]*(24)+in_buf[47]*(29)+in_buf[48]*(29)+in_buf[49]*(21)+in_buf[50]*(20)+in_buf[51]*(12)+in_buf[52]*(0)+in_buf[53]*(3)+in_buf[54]*(3)+in_buf[55]*(-2)+in_buf[56]*(2)+in_buf[57]*(0)+in_buf[58]*(17)+in_buf[59]*(23)+in_buf[60]*(40)+in_buf[61]*(4)+in_buf[62]*(15)+in_buf[63]*(13)+in_buf[64]*(13)+in_buf[65]*(-8)+in_buf[66]*(3)+in_buf[67]*(16)+in_buf[68]*(4)+in_buf[69]*(-3)+in_buf[70]*(2)+in_buf[71]*(19)+in_buf[72]*(16)+in_buf[73]*(14)+in_buf[74]*(23)+in_buf[75]*(20)+in_buf[76]*(20)+in_buf[77]*(19)+in_buf[78]*(37)+in_buf[79]*(30)+in_buf[80]*(-8)+in_buf[81]*(-5)+in_buf[82]*(1)+in_buf[83]*(3)+in_buf[84]*(-2)+in_buf[85]*(-1)+in_buf[86]*(-10)+in_buf[87]*(32)+in_buf[88]*(33)+in_buf[89]*(43)+in_buf[90]*(48)+in_buf[91]*(34)+in_buf[92]*(48)+in_buf[93]*(34)+in_buf[94]*(13)+in_buf[95]*(9)+in_buf[96]*(11)+in_buf[97]*(10)+in_buf[98]*(-2)+in_buf[99]*(5)+in_buf[100]*(2)+in_buf[101]*(8)+in_buf[102]*(12)+in_buf[103]*(17)+in_buf[104]*(13)+in_buf[105]*(23)+in_buf[106]*(23)+in_buf[107]*(27)+in_buf[108]*(23)+in_buf[109]*(-20)+in_buf[110]*(13)+in_buf[111]*(-1)+in_buf[112]*(-2)+in_buf[113]*(0)+in_buf[114]*(5)+in_buf[115]*(11)+in_buf[116]*(40)+in_buf[117]*(35)+in_buf[118]*(25)+in_buf[119]*(25)+in_buf[120]*(32)+in_buf[121]*(14)+in_buf[122]*(8)+in_buf[123]*(8)+in_buf[124]*(-10)+in_buf[125]*(-4)+in_buf[126]*(1)+in_buf[127]*(-8)+in_buf[128]*(-4)+in_buf[129]*(10)+in_buf[130]*(17)+in_buf[131]*(18)+in_buf[132]*(18)+in_buf[133]*(-3)+in_buf[134]*(-10)+in_buf[135]*(9)+in_buf[136]*(-12)+in_buf[137]*(-11)+in_buf[138]*(15)+in_buf[139]*(18)+in_buf[140]*(3)+in_buf[141]*(0)+in_buf[142]*(47)+in_buf[143]*(21)+in_buf[144]*(36)+in_buf[145]*(6)+in_buf[146]*(-1)+in_buf[147]*(2)+in_buf[148]*(-7)+in_buf[149]*(-10)+in_buf[150]*(-12)+in_buf[151]*(-17)+in_buf[152]*(-17)+in_buf[153]*(-5)+in_buf[154]*(-14)+in_buf[155]*(-11)+in_buf[156]*(2)+in_buf[157]*(1)+in_buf[158]*(-1)+in_buf[159]*(8)+in_buf[160]*(21)+in_buf[161]*(11)+in_buf[162]*(-1)+in_buf[163]*(3)+in_buf[164]*(0)+in_buf[165]*(-2)+in_buf[166]*(45)+in_buf[167]*(27)+in_buf[168]*(2)+in_buf[169]*(23)+in_buf[170]*(-13)+in_buf[171]*(6)+in_buf[172]*(40)+in_buf[173]*(19)+in_buf[174]*(0)+in_buf[175]*(-4)+in_buf[176]*(-4)+in_buf[177]*(-14)+in_buf[178]*(-25)+in_buf[179]*(-19)+in_buf[180]*(-22)+in_buf[181]*(-19)+in_buf[182]*(-10)+in_buf[183]*(-9)+in_buf[184]*(-13)+in_buf[185]*(-18)+in_buf[186]*(-18)+in_buf[187]*(-17)+in_buf[188]*(-9)+in_buf[189]*(-14)+in_buf[190]*(-7)+in_buf[191]*(-12)+in_buf[192]*(17)+in_buf[193]*(25)+in_buf[194]*(7)+in_buf[195]*(23)+in_buf[196]*(-1)+in_buf[197]*(28)+in_buf[198]*(-31)+in_buf[199]*(9)+in_buf[200]*(47)+in_buf[201]*(20)+in_buf[202]*(-12)+in_buf[203]*(0)+in_buf[204]*(6)+in_buf[205]*(-4)+in_buf[206]*(-17)+in_buf[207]*(-12)+in_buf[208]*(-11)+in_buf[209]*(-18)+in_buf[210]*(-6)+in_buf[211]*(-8)+in_buf[212]*(-21)+in_buf[213]*(-27)+in_buf[214]*(-17)+in_buf[215]*(-21)+in_buf[216]*(-19)+in_buf[217]*(-29)+in_buf[218]*(-33)+in_buf[219]*(-27)+in_buf[220]*(5)+in_buf[221]*(4)+in_buf[222]*(2)+in_buf[223]*(19)+in_buf[224]*(23)+in_buf[225]*(18)+in_buf[226]*(-48)+in_buf[227]*(10)+in_buf[228]*(30)+in_buf[229]*(19)+in_buf[230]*(-8)+in_buf[231]*(7)+in_buf[232]*(9)+in_buf[233]*(-9)+in_buf[234]*(-13)+in_buf[235]*(-18)+in_buf[236]*(-20)+in_buf[237]*(-22)+in_buf[238]*(-12)+in_buf[239]*(-28)+in_buf[240]*(-32)+in_buf[241]*(-26)+in_buf[242]*(-37)+in_buf[243]*(-17)+in_buf[244]*(-4)+in_buf[245]*(-17)+in_buf[246]*(-4)+in_buf[247]*(-30)+in_buf[248]*(-40)+in_buf[249]*(-38)+in_buf[250]*(-26)+in_buf[251]*(-6)+in_buf[252]*(3)+in_buf[253]*(-20)+in_buf[254]*(-36)+in_buf[255]*(3)+in_buf[256]*(15)+in_buf[257]*(1)+in_buf[258]*(-14)+in_buf[259]*(6)+in_buf[260]*(11)+in_buf[261]*(-15)+in_buf[262]*(-29)+in_buf[263]*(-21)+in_buf[264]*(-22)+in_buf[265]*(-12)+in_buf[266]*(-5)+in_buf[267]*(-24)+in_buf[268]*(-12)+in_buf[269]*(-15)+in_buf[270]*(-19)+in_buf[271]*(-21)+in_buf[272]*(-3)+in_buf[273]*(1)+in_buf[274]*(13)+in_buf[275]*(-8)+in_buf[276]*(-29)+in_buf[277]*(-33)+in_buf[278]*(-33)+in_buf[279]*(-22)+in_buf[280]*(5)+in_buf[281]*(-6)+in_buf[282]*(7)+in_buf[283]*(-19)+in_buf[284]*(-4)+in_buf[285]*(-10)+in_buf[286]*(-10)+in_buf[287]*(-1)+in_buf[288]*(9)+in_buf[289]*(-7)+in_buf[290]*(-9)+in_buf[291]*(-10)+in_buf[292]*(4)+in_buf[293]*(10)+in_buf[294]*(10)+in_buf[295]*(3)+in_buf[296]*(2)+in_buf[297]*(0)+in_buf[298]*(-4)+in_buf[299]*(-11)+in_buf[300]*(-15)+in_buf[301]*(0)+in_buf[302]*(-2)+in_buf[303]*(0)+in_buf[304]*(0)+in_buf[305]*(-39)+in_buf[306]*(-24)+in_buf[307]*(-38)+in_buf[308]*(1)+in_buf[309]*(-21)+in_buf[310]*(7)+in_buf[311]*(-10)+in_buf[312]*(-6)+in_buf[313]*(4)+in_buf[314]*(0)+in_buf[315]*(16)+in_buf[316]*(9)+in_buf[317]*(18)+in_buf[318]*(6)+in_buf[319]*(8)+in_buf[320]*(12)+in_buf[321]*(16)+in_buf[322]*(28)+in_buf[323]*(15)+in_buf[324]*(11)+in_buf[325]*(14)+in_buf[326]*(18)+in_buf[327]*(-2)+in_buf[328]*(6)+in_buf[329]*(7)+in_buf[330]*(11)+in_buf[331]*(8)+in_buf[332]*(10)+in_buf[333]*(-28)+in_buf[334]*(0)+in_buf[335]*(-10)+in_buf[336]*(2)+in_buf[337]*(-18)+in_buf[338]*(-22)+in_buf[339]*(-9)+in_buf[340]*(0)+in_buf[341]*(15)+in_buf[342]*(15)+in_buf[343]*(31)+in_buf[344]*(29)+in_buf[345]*(36)+in_buf[346]*(22)+in_buf[347]*(12)+in_buf[348]*(0)+in_buf[349]*(14)+in_buf[350]*(34)+in_buf[351]*(22)+in_buf[352]*(18)+in_buf[353]*(27)+in_buf[354]*(16)+in_buf[355]*(11)+in_buf[356]*(17)+in_buf[357]*(1)+in_buf[358]*(16)+in_buf[359]*(27)+in_buf[360]*(22)+in_buf[361]*(12)+in_buf[362]*(18)+in_buf[363]*(-8)+in_buf[364]*(24)+in_buf[365]*(-6)+in_buf[366]*(-5)+in_buf[367]*(19)+in_buf[368]*(-9)+in_buf[369]*(25)+in_buf[370]*(22)+in_buf[371]*(6)+in_buf[372]*(7)+in_buf[373]*(13)+in_buf[374]*(10)+in_buf[375]*(-6)+in_buf[376]*(-6)+in_buf[377]*(-1)+in_buf[378]*(24)+in_buf[379]*(29)+in_buf[380]*(20)+in_buf[381]*(8)+in_buf[382]*(16)+in_buf[383]*(20)+in_buf[384]*(1)+in_buf[385]*(4)+in_buf[386]*(-2)+in_buf[387]*(30)+in_buf[388]*(17)+in_buf[389]*(9)+in_buf[390]*(2)+in_buf[391]*(-11)+in_buf[392]*(17)+in_buf[393]*(10)+in_buf[394]*(32)+in_buf[395]*(37)+in_buf[396]*(-23)+in_buf[397]*(15)+in_buf[398]*(-4)+in_buf[399]*(-26)+in_buf[400]*(-14)+in_buf[401]*(-3)+in_buf[402]*(0)+in_buf[403]*(-11)+in_buf[404]*(-16)+in_buf[405]*(2)+in_buf[406]*(18)+in_buf[407]*(14)+in_buf[408]*(6)+in_buf[409]*(2)+in_buf[410]*(26)+in_buf[411]*(19)+in_buf[412]*(13)+in_buf[413]*(10)+in_buf[414]*(6)+in_buf[415]*(3)+in_buf[416]*(-10)+in_buf[417]*(-19)+in_buf[418]*(-27)+in_buf[419]*(-7)+in_buf[420]*(12)+in_buf[421]*(17)+in_buf[422]*(37)+in_buf[423]*(0)+in_buf[424]*(-13)+in_buf[425]*(-4)+in_buf[426]*(-9)+in_buf[427]*(-23)+in_buf[428]*(-18)+in_buf[429]*(-16)+in_buf[430]*(-33)+in_buf[431]*(-41)+in_buf[432]*(-12)+in_buf[433]*(8)+in_buf[434]*(15)+in_buf[435]*(-6)+in_buf[436]*(-5)+in_buf[437]*(-2)+in_buf[438]*(20)+in_buf[439]*(15)+in_buf[440]*(15)+in_buf[441]*(21)+in_buf[442]*(-6)+in_buf[443]*(-15)+in_buf[444]*(-15)+in_buf[445]*(-25)+in_buf[446]*(-42)+in_buf[447]*(-18)+in_buf[448]*(-1)+in_buf[449]*(17)+in_buf[450]*(33)+in_buf[451]*(15)+in_buf[452]*(-10)+in_buf[453]*(-9)+in_buf[454]*(-27)+in_buf[455]*(-12)+in_buf[456]*(-22)+in_buf[457]*(-5)+in_buf[458]*(-12)+in_buf[459]*(-6)+in_buf[460]*(0)+in_buf[461]*(13)+in_buf[462]*(15)+in_buf[463]*(-11)+in_buf[464]*(-19)+in_buf[465]*(-9)+in_buf[466]*(29)+in_buf[467]*(16)+in_buf[468]*(11)+in_buf[469]*(5)+in_buf[470]*(-3)+in_buf[471]*(-7)+in_buf[472]*(-9)+in_buf[473]*(-24)+in_buf[474]*(-45)+in_buf[475]*(-16)+in_buf[476]*(2)+in_buf[477]*(16)+in_buf[478]*(21)+in_buf[479]*(26)+in_buf[480]*(2)+in_buf[481]*(-13)+in_buf[482]*(-14)+in_buf[483]*(1)+in_buf[484]*(-1)+in_buf[485]*(-15)+in_buf[486]*(-2)+in_buf[487]*(13)+in_buf[488]*(-4)+in_buf[489]*(9)+in_buf[490]*(3)+in_buf[491]*(-6)+in_buf[492]*(4)+in_buf[493]*(2)+in_buf[494]*(9)+in_buf[495]*(23)+in_buf[496]*(11)+in_buf[497]*(0)+in_buf[498]*(-15)+in_buf[499]*(-6)+in_buf[500]*(-20)+in_buf[501]*(-32)+in_buf[502]*(-48)+in_buf[503]*(-6)+in_buf[504]*(23)+in_buf[505]*(17)+in_buf[506]*(33)+in_buf[507]*(44)+in_buf[508]*(-4)+in_buf[509]*(1)+in_buf[510]*(3)+in_buf[511]*(26)+in_buf[512]*(21)+in_buf[513]*(12)+in_buf[514]*(14)+in_buf[515]*(8)+in_buf[516]*(8)+in_buf[517]*(10)+in_buf[518]*(4)+in_buf[519]*(18)+in_buf[520]*(11)+in_buf[521]*(9)+in_buf[522]*(15)+in_buf[523]*(3)+in_buf[524]*(-16)+in_buf[525]*(-26)+in_buf[526]*(-31)+in_buf[527]*(-16)+in_buf[528]*(-22)+in_buf[529]*(-2)+in_buf[530]*(-25)+in_buf[531]*(0)+in_buf[532]*(24)+in_buf[533]*(38)+in_buf[534]*(25)+in_buf[535]*(41)+in_buf[536]*(5)+in_buf[537]*(0)+in_buf[538]*(13)+in_buf[539]*(17)+in_buf[540]*(20)+in_buf[541]*(33)+in_buf[542]*(32)+in_buf[543]*(25)+in_buf[544]*(16)+in_buf[545]*(13)+in_buf[546]*(21)+in_buf[547]*(16)+in_buf[548]*(0)+in_buf[549]*(11)+in_buf[550]*(11)+in_buf[551]*(-7)+in_buf[552]*(-14)+in_buf[553]*(-26)+in_buf[554]*(-26)+in_buf[555]*(0)+in_buf[556]*(0)+in_buf[557]*(13)+in_buf[558]*(-19)+in_buf[559]*(2)+in_buf[560]*(0)+in_buf[561]*(-11)+in_buf[562]*(-3)+in_buf[563]*(16)+in_buf[564]*(6)+in_buf[565]*(-10)+in_buf[566]*(-11)+in_buf[567]*(17)+in_buf[568]*(22)+in_buf[569]*(36)+in_buf[570]*(33)+in_buf[571]*(11)+in_buf[572]*(11)+in_buf[573]*(17)+in_buf[574]*(27)+in_buf[575]*(14)+in_buf[576]*(-2)+in_buf[577]*(-6)+in_buf[578]*(0)+in_buf[579]*(-10)+in_buf[580]*(-16)+in_buf[581]*(-23)+in_buf[582]*(-14)+in_buf[583]*(-40)+in_buf[584]*(-31)+in_buf[585]*(-19)+in_buf[586]*(-1)+in_buf[587]*(8)+in_buf[588]*(2)+in_buf[589]*(4)+in_buf[590]*(-25)+in_buf[591]*(-2)+in_buf[592]*(-15)+in_buf[593]*(-40)+in_buf[594]*(-15)+in_buf[595]*(11)+in_buf[596]*(9)+in_buf[597]*(24)+in_buf[598]*(24)+in_buf[599]*(18)+in_buf[600]*(14)+in_buf[601]*(17)+in_buf[602]*(14)+in_buf[603]*(3)+in_buf[604]*(1)+in_buf[605]*(11)+in_buf[606]*(21)+in_buf[607]*(-2)+in_buf[608]*(-24)+in_buf[609]*(-27)+in_buf[610]*(-40)+in_buf[611]*(-51)+in_buf[612]*(-33)+in_buf[613]*(2)+in_buf[614]*(28)+in_buf[615]*(2)+in_buf[616]*(3)+in_buf[617]*(10)+in_buf[618]*(-3)+in_buf[619]*(-11)+in_buf[620]*(-16)+in_buf[621]*(-19)+in_buf[622]*(-12)+in_buf[623]*(-6)+in_buf[624]*(1)+in_buf[625]*(19)+in_buf[626]*(21)+in_buf[627]*(11)+in_buf[628]*(11)+in_buf[629]*(12)+in_buf[630]*(-2)+in_buf[631]*(6)+in_buf[632]*(6)+in_buf[633]*(3)+in_buf[634]*(-16)+in_buf[635]*(-16)+in_buf[636]*(-25)+in_buf[637]*(-60)+in_buf[638]*(-47)+in_buf[639]*(-50)+in_buf[640]*(-30)+in_buf[641]*(4)+in_buf[642]*(35)+in_buf[643]*(0)+in_buf[644]*(2)+in_buf[645]*(0)+in_buf[646]*(27)+in_buf[647]*(12)+in_buf[648]*(10)+in_buf[649]*(-4)+in_buf[650]*(-20)+in_buf[651]*(-32)+in_buf[652]*(-25)+in_buf[653]*(0)+in_buf[654]*(-5)+in_buf[655]*(-1)+in_buf[656]*(6)+in_buf[657]*(-4)+in_buf[658]*(-12)+in_buf[659]*(-19)+in_buf[660]*(-35)+in_buf[661]*(-48)+in_buf[662]*(-60)+in_buf[663]*(-34)+in_buf[664]*(-18)+in_buf[665]*(-22)+in_buf[666]*(-46)+in_buf[667]*(-40)+in_buf[668]*(-32)+in_buf[669]*(-17)+in_buf[670]*(13)+in_buf[671]*(-2)+in_buf[672]*(4)+in_buf[673]*(1)+in_buf[674]*(0)+in_buf[675]*(31)+in_buf[676]*(-11)+in_buf[677]*(-8)+in_buf[678]*(-21)+in_buf[679]*(-48)+in_buf[680]*(-45)+in_buf[681]*(-31)+in_buf[682]*(-22)+in_buf[683]*(-12)+in_buf[684]*(-13)+in_buf[685]*(-27)+in_buf[686]*(-8)+in_buf[687]*(-29)+in_buf[688]*(-34)+in_buf[689]*(-54)+in_buf[690]*(-52)+in_buf[691]*(-20)+in_buf[692]*(6)+in_buf[693]*(10)+in_buf[694]*(-28)+in_buf[695]*(-37)+in_buf[696]*(-17)+in_buf[697]*(20)+in_buf[698]*(9)+in_buf[699]*(4)+in_buf[700]*(2)+in_buf[701]*(2)+in_buf[702]*(-1)+in_buf[703]*(1)+in_buf[704]*(-3)+in_buf[705]*(-5)+in_buf[706]*(1)+in_buf[707]*(-29)+in_buf[708]*(-51)+in_buf[709]*(-45)+in_buf[710]*(-51)+in_buf[711]*(-60)+in_buf[712]*(-27)+in_buf[713]*(-40)+in_buf[714]*(-45)+in_buf[715]*(-49)+in_buf[716]*(-22)+in_buf[717]*(-22)+in_buf[718]*(-21)+in_buf[719]*(4)+in_buf[720]*(11)+in_buf[721]*(7)+in_buf[722]*(15)+in_buf[723]*(-22)+in_buf[724]*(-30)+in_buf[725]*(-1)+in_buf[726]*(2)+in_buf[727]*(2)+in_buf[728]*(4)+in_buf[729]*(2)+in_buf[730]*(-1)+in_buf[731]*(-6)+in_buf[732]*(6)+in_buf[733]*(34)+in_buf[734]*(14)+in_buf[735]*(-8)+in_buf[736]*(-16)+in_buf[737]*(-34)+in_buf[738]*(-32)+in_buf[739]*(-27)+in_buf[740]*(-52)+in_buf[741]*(-47)+in_buf[742]*(-69)+in_buf[743]*(-41)+in_buf[744]*(-5)+in_buf[745]*(-23)+in_buf[746]*(-55)+in_buf[747]*(-3)+in_buf[748]*(17)+in_buf[749]*(3)+in_buf[750]*(-3)+in_buf[751]*(-22)+in_buf[752]*(0)+in_buf[753]*(1)+in_buf[754]*(-1)+in_buf[755]*(3)+in_buf[756]*(-3)+in_buf[757]*(-1)+in_buf[758]*(-3)+in_buf[759]*(-3)+in_buf[760]*(11)+in_buf[761]*(1)+in_buf[762]*(6)+in_buf[763]*(10)+in_buf[764]*(9)+in_buf[765]*(13)+in_buf[766]*(-23)+in_buf[767]*(0)+in_buf[768]*(3)+in_buf[769]*(-2)+in_buf[770]*(-29)+in_buf[771]*(-33)+in_buf[772]*(6)+in_buf[773]*(-21)+in_buf[774]*(-22)+in_buf[775]*(-17)+in_buf[776]*(17)+in_buf[777]*(15)+in_buf[778]*(14)+in_buf[779]*(0)+in_buf[780]*(0)+in_buf[781]*(-2)+in_buf[782]*(0)+in_buf[783]*(4);
assign in_buf_weight04=in_buf[0]*(1)+in_buf[1]*(2)+in_buf[2]*(0)+in_buf[3]*(-2)+in_buf[4]*(4)+in_buf[5]*(-1)+in_buf[6]*(0)+in_buf[7]*(1)+in_buf[8]*(3)+in_buf[9]*(4)+in_buf[10]*(-1)+in_buf[11]*(0)+in_buf[12]*(0)+in_buf[13]*(-3)+in_buf[14]*(5)+in_buf[15]*(3)+in_buf[16]*(-1)+in_buf[17]*(-1)+in_buf[18]*(-3)+in_buf[19]*(0)+in_buf[20]*(2)+in_buf[21]*(-3)+in_buf[22]*(1)+in_buf[23]*(-3)+in_buf[24]*(0)+in_buf[25]*(2)+in_buf[26]*(-3)+in_buf[27]*(-1)+in_buf[28]*(0)+in_buf[29]*(4)+in_buf[30]*(1)+in_buf[31]*(4)+in_buf[32]*(-6)+in_buf[33]*(-6)+in_buf[34]*(-1)+in_buf[35]*(-9)+in_buf[36]*(-3)+in_buf[37]*(-1)+in_buf[38]*(-10)+in_buf[39]*(-14)+in_buf[40]*(-26)+in_buf[41]*(-34)+in_buf[42]*(-7)+in_buf[43]*(-6)+in_buf[44]*(-12)+in_buf[45]*(-17)+in_buf[46]*(-20)+in_buf[47]*(-21)+in_buf[48]*(-15)+in_buf[49]*(-11)+in_buf[50]*(-12)+in_buf[51]*(-15)+in_buf[52]*(4)+in_buf[53]*(-2)+in_buf[54]*(2)+in_buf[55]*(5)+in_buf[56]*(-1)+in_buf[57]*(-2)+in_buf[58]*(-12)+in_buf[59]*(-24)+in_buf[60]*(-32)+in_buf[61]*(-12)+in_buf[62]*(-6)+in_buf[63]*(-4)+in_buf[64]*(-22)+in_buf[65]*(-12)+in_buf[66]*(-11)+in_buf[67]*(-20)+in_buf[68]*(-37)+in_buf[69]*(-24)+in_buf[70]*(-9)+in_buf[71]*(2)+in_buf[72]*(-31)+in_buf[73]*(-13)+in_buf[74]*(21)+in_buf[75]*(1)+in_buf[76]*(3)+in_buf[77]*(-7)+in_buf[78]*(-5)+in_buf[79]*(-10)+in_buf[80]*(4)+in_buf[81]*(9)+in_buf[82]*(0)+in_buf[83]*(-1)+in_buf[84]*(1)+in_buf[85]*(3)+in_buf[86]*(6)+in_buf[87]*(-27)+in_buf[88]*(-29)+in_buf[89]*(-12)+in_buf[90]*(-18)+in_buf[91]*(-40)+in_buf[92]*(-43)+in_buf[93]*(-43)+in_buf[94]*(-30)+in_buf[95]*(-25)+in_buf[96]*(-31)+in_buf[97]*(-19)+in_buf[98]*(-22)+in_buf[99]*(0)+in_buf[100]*(6)+in_buf[101]*(-18)+in_buf[102]*(-29)+in_buf[103]*(-42)+in_buf[104]*(-17)+in_buf[105]*(9)+in_buf[106]*(-2)+in_buf[107]*(7)+in_buf[108]*(0)+in_buf[109]*(20)+in_buf[110]*(-6)+in_buf[111]*(1)+in_buf[112]*(-3)+in_buf[113]*(0)+in_buf[114]*(-4)+in_buf[115]*(-27)+in_buf[116]*(-34)+in_buf[117]*(-35)+in_buf[118]*(-33)+in_buf[119]*(-7)+in_buf[120]*(-18)+in_buf[121]*(-18)+in_buf[122]*(0)+in_buf[123]*(7)+in_buf[124]*(8)+in_buf[125]*(0)+in_buf[126]*(0)+in_buf[127]*(4)+in_buf[128]*(13)+in_buf[129]*(-1)+in_buf[130]*(-10)+in_buf[131]*(-21)+in_buf[132]*(-13)+in_buf[133]*(7)+in_buf[134]*(-8)+in_buf[135]*(6)+in_buf[136]*(48)+in_buf[137]*(34)+in_buf[138]*(41)+in_buf[139]*(7)+in_buf[140]*(3)+in_buf[141]*(0)+in_buf[142]*(-15)+in_buf[143]*(-16)+in_buf[144]*(-32)+in_buf[145]*(-50)+in_buf[146]*(-15)+in_buf[147]*(-8)+in_buf[148]*(-27)+in_buf[149]*(-1)+in_buf[150]*(-2)+in_buf[151]*(12)+in_buf[152]*(17)+in_buf[153]*(4)+in_buf[154]*(2)+in_buf[155]*(-3)+in_buf[156]*(-5)+in_buf[157]*(-2)+in_buf[158]*(-6)+in_buf[159]*(2)+in_buf[160]*(9)+in_buf[161]*(10)+in_buf[162]*(8)+in_buf[163]*(9)+in_buf[164]*(27)+in_buf[165]*(44)+in_buf[166]*(17)+in_buf[167]*(-7)+in_buf[168]*(0)+in_buf[169]*(-17)+in_buf[170]*(-12)+in_buf[171]*(-42)+in_buf[172]*(-66)+in_buf[173]*(-52)+in_buf[174]*(-26)+in_buf[175]*(-11)+in_buf[176]*(-3)+in_buf[177]*(3)+in_buf[178]*(-1)+in_buf[179]*(2)+in_buf[180]*(5)+in_buf[181]*(6)+in_buf[182]*(5)+in_buf[183]*(0)+in_buf[184]*(-2)+in_buf[185]*(0)+in_buf[186]*(-11)+in_buf[187]*(8)+in_buf[188]*(10)+in_buf[189]*(13)+in_buf[190]*(17)+in_buf[191]*(24)+in_buf[192]*(12)+in_buf[193]*(44)+in_buf[194]*(7)+in_buf[195]*(-15)+in_buf[196]*(2)+in_buf[197]*(-31)+in_buf[198]*(-29)+in_buf[199]*(-57)+in_buf[200]*(-34)+in_buf[201]*(-47)+in_buf[202]*(-12)+in_buf[203]*(-13)+in_buf[204]*(17)+in_buf[205]*(0)+in_buf[206]*(-3)+in_buf[207]*(-4)+in_buf[208]*(5)+in_buf[209]*(7)+in_buf[210]*(0)+in_buf[211]*(10)+in_buf[212]*(0)+in_buf[213]*(-15)+in_buf[214]*(-13)+in_buf[215]*(0)+in_buf[216]*(9)+in_buf[217]*(13)+in_buf[218]*(18)+in_buf[219]*(16)+in_buf[220]*(26)+in_buf[221]*(41)+in_buf[222]*(-7)+in_buf[223]*(-22)+in_buf[224]*(-17)+in_buf[225]*(-19)+in_buf[226]*(-20)+in_buf[227]*(3)+in_buf[228]*(-20)+in_buf[229]*(-9)+in_buf[230]*(0)+in_buf[231]*(7)+in_buf[232]*(10)+in_buf[233]*(-6)+in_buf[234]*(0)+in_buf[235]*(6)+in_buf[236]*(15)+in_buf[237]*(20)+in_buf[238]*(15)+in_buf[239]*(3)+in_buf[240]*(0)+in_buf[241]*(-11)+in_buf[242]*(0)+in_buf[243]*(2)+in_buf[244]*(2)+in_buf[245]*(13)+in_buf[246]*(2)+in_buf[247]*(4)+in_buf[248]*(32)+in_buf[249]*(35)+in_buf[250]*(36)+in_buf[251]*(17)+in_buf[252]*(-8)+in_buf[253]*(-25)+in_buf[254]*(-4)+in_buf[255]*(19)+in_buf[256]*(-22)+in_buf[257]*(3)+in_buf[258]*(13)+in_buf[259]*(-1)+in_buf[260]*(1)+in_buf[261]*(7)+in_buf[262]*(16)+in_buf[263]*(17)+in_buf[264]*(17)+in_buf[265]*(31)+in_buf[266]*(18)+in_buf[267]*(0)+in_buf[268]*(-5)+in_buf[269]*(-3)+in_buf[270]*(-14)+in_buf[271]*(-11)+in_buf[272]*(0)+in_buf[273]*(4)+in_buf[274]*(8)+in_buf[275]*(14)+in_buf[276]*(9)+in_buf[277]*(36)+in_buf[278]*(28)+in_buf[279]*(-10)+in_buf[280]*(-14)+in_buf[281]*(-12)+in_buf[282]*(-32)+in_buf[283]*(2)+in_buf[284]*(15)+in_buf[285]*(19)+in_buf[286]*(19)+in_buf[287]*(-2)+in_buf[288]*(-3)+in_buf[289]*(4)+in_buf[290]*(21)+in_buf[291]*(21)+in_buf[292]*(32)+in_buf[293]*(15)+in_buf[294]*(9)+in_buf[295]*(-10)+in_buf[296]*(-21)+in_buf[297]*(-31)+in_buf[298]*(-29)+in_buf[299]*(-12)+in_buf[300]*(5)+in_buf[301]*(8)+in_buf[302]*(-3)+in_buf[303]*(16)+in_buf[304]*(-2)+in_buf[305]*(1)+in_buf[306]*(6)+in_buf[307]*(13)+in_buf[308]*(-18)+in_buf[309]*(-37)+in_buf[310]*(-24)+in_buf[311]*(0)+in_buf[312]*(31)+in_buf[313]*(38)+in_buf[314]*(16)+in_buf[315]*(7)+in_buf[316]*(9)+in_buf[317]*(21)+in_buf[318]*(16)+in_buf[319]*(7)+in_buf[320]*(21)+in_buf[321]*(10)+in_buf[322]*(12)+in_buf[323]*(-11)+in_buf[324]*(-24)+in_buf[325]*(-30)+in_buf[326]*(-26)+in_buf[327]*(-6)+in_buf[328]*(14)+in_buf[329]*(4)+in_buf[330]*(0)+in_buf[331]*(-4)+in_buf[332]*(-2)+in_buf[333]*(4)+in_buf[334]*(30)+in_buf[335]*(-21)+in_buf[336]*(-12)+in_buf[337]*(-16)+in_buf[338]*(-11)+in_buf[339]*(22)+in_buf[340]*(45)+in_buf[341]*(38)+in_buf[342]*(23)+in_buf[343]*(19)+in_buf[344]*(10)+in_buf[345]*(7)+in_buf[346]*(-3)+in_buf[347]*(-6)+in_buf[348]*(-12)+in_buf[349]*(4)+in_buf[350]*(-10)+in_buf[351]*(-13)+in_buf[352]*(-9)+in_buf[353]*(4)+in_buf[354]*(-8)+in_buf[355]*(16)+in_buf[356]*(22)+in_buf[357]*(15)+in_buf[358]*(2)+in_buf[359]*(-9)+in_buf[360]*(-13)+in_buf[361]*(-13)+in_buf[362]*(13)+in_buf[363]*(-20)+in_buf[364]*(10)+in_buf[365]*(-2)+in_buf[366]*(-24)+in_buf[367]*(10)+in_buf[368]*(13)+in_buf[369]*(21)+in_buf[370]*(7)+in_buf[371]*(20)+in_buf[372]*(7)+in_buf[373]*(3)+in_buf[374]*(-16)+in_buf[375]*(-7)+in_buf[376]*(-2)+in_buf[377]*(11)+in_buf[378]*(11)+in_buf[379]*(6)+in_buf[380]*(1)+in_buf[381]*(6)+in_buf[382]*(-3)+in_buf[383]*(9)+in_buf[384]*(20)+in_buf[385]*(5)+in_buf[386]*(6)+in_buf[387]*(-20)+in_buf[388]*(-39)+in_buf[389]*(-4)+in_buf[390]*(26)+in_buf[391]*(38)+in_buf[392]*(-3)+in_buf[393]*(-4)+in_buf[394]*(-14)+in_buf[395]*(18)+in_buf[396]*(-7)+in_buf[397]*(4)+in_buf[398]*(13)+in_buf[399]*(0)+in_buf[400]*(2)+in_buf[401]*(-11)+in_buf[402]*(-10)+in_buf[403]*(-5)+in_buf[404]*(-1)+in_buf[405]*(15)+in_buf[406]*(12)+in_buf[407]*(7)+in_buf[408]*(17)+in_buf[409]*(0)+in_buf[410]*(-19)+in_buf[411]*(-2)+in_buf[412]*(3)+in_buf[413]*(-9)+in_buf[414]*(-9)+in_buf[415]*(-28)+in_buf[416]*(-29)+in_buf[417]*(-10)+in_buf[418]*(45)+in_buf[419]*(15)+in_buf[420]*(-9)+in_buf[421]*(-3)+in_buf[422]*(-27)+in_buf[423]*(14)+in_buf[424]*(-16)+in_buf[425]*(0)+in_buf[426]*(8)+in_buf[427]*(-15)+in_buf[428]*(-10)+in_buf[429]*(-11)+in_buf[430]*(-8)+in_buf[431]*(3)+in_buf[432]*(3)+in_buf[433]*(19)+in_buf[434]*(24)+in_buf[435]*(16)+in_buf[436]*(11)+in_buf[437]*(-3)+in_buf[438]*(-7)+in_buf[439]*(0)+in_buf[440]*(-9)+in_buf[441]*(-27)+in_buf[442]*(-21)+in_buf[443]*(-37)+in_buf[444]*(-28)+in_buf[445]*(-7)+in_buf[446]*(33)+in_buf[447]*(8)+in_buf[448]*(2)+in_buf[449]*(-3)+in_buf[450]*(-20)+in_buf[451]*(-4)+in_buf[452]*(-12)+in_buf[453]*(-10)+in_buf[454]*(10)+in_buf[455]*(-10)+in_buf[456]*(-22)+in_buf[457]*(-17)+in_buf[458]*(-1)+in_buf[459]*(4)+in_buf[460]*(16)+in_buf[461]*(18)+in_buf[462]*(23)+in_buf[463]*(14)+in_buf[464]*(14)+in_buf[465]*(1)+in_buf[466]*(-3)+in_buf[467]*(-22)+in_buf[468]*(-18)+in_buf[469]*(-15)+in_buf[470]*(-18)+in_buf[471]*(-30)+in_buf[472]*(-17)+in_buf[473]*(0)+in_buf[474]*(34)+in_buf[475]*(4)+in_buf[476]*(2)+in_buf[477]*(-5)+in_buf[478]*(-27)+in_buf[479]*(2)+in_buf[480]*(-14)+in_buf[481]*(-9)+in_buf[482]*(0)+in_buf[483]*(-14)+in_buf[484]*(-7)+in_buf[485]*(-11)+in_buf[486]*(0)+in_buf[487]*(10)+in_buf[488]*(17)+in_buf[489]*(19)+in_buf[490]*(5)+in_buf[491]*(0)+in_buf[492]*(9)+in_buf[493]*(-1)+in_buf[494]*(0)+in_buf[495]*(-16)+in_buf[496]*(-5)+in_buf[497]*(3)+in_buf[498]*(-17)+in_buf[499]*(-13)+in_buf[500]*(5)+in_buf[501]*(-11)+in_buf[502]*(13)+in_buf[503]*(25)+in_buf[504]*(-3)+in_buf[505]*(-7)+in_buf[506]*(-22)+in_buf[507]*(3)+in_buf[508]*(0)+in_buf[509]*(-2)+in_buf[510]*(13)+in_buf[511]*(-7)+in_buf[512]*(0)+in_buf[513]*(-8)+in_buf[514]*(0)+in_buf[515]*(9)+in_buf[516]*(5)+in_buf[517]*(9)+in_buf[518]*(4)+in_buf[519]*(0)+in_buf[520]*(-13)+in_buf[521]*(-4)+in_buf[522]*(-12)+in_buf[523]*(-3)+in_buf[524]*(16)+in_buf[525]*(0)+in_buf[526]*(3)+in_buf[527]*(0)+in_buf[528]*(5)+in_buf[529]*(0)+in_buf[530]*(-10)+in_buf[531]*(23)+in_buf[532]*(10)+in_buf[533]*(-35)+in_buf[534]*(-12)+in_buf[535]*(-30)+in_buf[536]*(-12)+in_buf[537]*(-7)+in_buf[538]*(-4)+in_buf[539]*(-2)+in_buf[540]*(5)+in_buf[541]*(-1)+in_buf[542]*(5)+in_buf[543]*(-12)+in_buf[544]*(-21)+in_buf[545]*(-8)+in_buf[546]*(-7)+in_buf[547]*(0)+in_buf[548]*(-1)+in_buf[549]*(-5)+in_buf[550]*(-5)+in_buf[551]*(4)+in_buf[552]*(0)+in_buf[553]*(1)+in_buf[554]*(11)+in_buf[555]*(35)+in_buf[556]*(21)+in_buf[557]*(26)+in_buf[558]*(26)+in_buf[559]*(-9)+in_buf[560]*(4)+in_buf[561]*(-4)+in_buf[562]*(-18)+in_buf[563]*(-22)+in_buf[564]*(-15)+in_buf[565]*(0)+in_buf[566]*(-5)+in_buf[567]*(-1)+in_buf[568]*(5)+in_buf[569]*(-3)+in_buf[570]*(8)+in_buf[571]*(-2)+in_buf[572]*(-21)+in_buf[573]*(-10)+in_buf[574]*(-7)+in_buf[575]*(-6)+in_buf[576]*(1)+in_buf[577]*(-1)+in_buf[578]*(-6)+in_buf[579]*(-5)+in_buf[580]*(8)+in_buf[581]*(10)+in_buf[582]*(21)+in_buf[583]*(33)+in_buf[584]*(31)+in_buf[585]*(34)+in_buf[586]*(0)+in_buf[587]*(5)+in_buf[588]*(-3)+in_buf[589]*(1)+in_buf[590]*(-15)+in_buf[591]*(-11)+in_buf[592]*(3)+in_buf[593]*(7)+in_buf[594]*(1)+in_buf[595]*(0)+in_buf[596]*(2)+in_buf[597]*(1)+in_buf[598]*(0)+in_buf[599]*(8)+in_buf[600]*(-2)+in_buf[601]*(-4)+in_buf[602]*(-7)+in_buf[603]*(-3)+in_buf[604]*(-4)+in_buf[605]*(2)+in_buf[606]*(-6)+in_buf[607]*(5)+in_buf[608]*(12)+in_buf[609]*(19)+in_buf[610]*(21)+in_buf[611]*(33)+in_buf[612]*(8)+in_buf[613]*(3)+in_buf[614]*(-20)+in_buf[615]*(-1)+in_buf[616]*(-8)+in_buf[617]*(-2)+in_buf[618]*(-18)+in_buf[619]*(-9)+in_buf[620]*(26)+in_buf[621]*(1)+in_buf[622]*(6)+in_buf[623]*(-2)+in_buf[624]*(0)+in_buf[625]*(6)+in_buf[626]*(-6)+in_buf[627]*(11)+in_buf[628]*(-1)+in_buf[629]*(-9)+in_buf[630]*(-5)+in_buf[631]*(-16)+in_buf[632]*(-8)+in_buf[633]*(-2)+in_buf[634]*(-2)+in_buf[635]*(-2)+in_buf[636]*(18)+in_buf[637]*(11)+in_buf[638]*(21)+in_buf[639]*(32)+in_buf[640]*(38)+in_buf[641]*(23)+in_buf[642]*(-10)+in_buf[643]*(-3)+in_buf[644]*(-3)+in_buf[645]*(0)+in_buf[646]*(-20)+in_buf[647]*(-18)+in_buf[648]*(28)+in_buf[649]*(0)+in_buf[650]*(-13)+in_buf[651]*(-17)+in_buf[652]*(-9)+in_buf[653]*(-4)+in_buf[654]*(-5)+in_buf[655]*(-11)+in_buf[656]*(-8)+in_buf[657]*(-3)+in_buf[658]*(-17)+in_buf[659]*(-2)+in_buf[660]*(4)+in_buf[661]*(5)+in_buf[662]*(13)+in_buf[663]*(12)+in_buf[664]*(18)+in_buf[665]*(8)+in_buf[666]*(28)+in_buf[667]*(50)+in_buf[668]*(25)+in_buf[669]*(13)+in_buf[670]*(-23)+in_buf[671]*(3)+in_buf[672]*(-2)+in_buf[673]*(0)+in_buf[674]*(-7)+in_buf[675]*(-29)+in_buf[676]*(-18)+in_buf[677]*(-15)+in_buf[678]*(0)+in_buf[679]*(-1)+in_buf[680]*(-2)+in_buf[681]*(-15)+in_buf[682]*(-2)+in_buf[683]*(-7)+in_buf[684]*(-9)+in_buf[685]*(0)+in_buf[686]*(-9)+in_buf[687]*(-4)+in_buf[688]*(2)+in_buf[689]*(-13)+in_buf[690]*(7)+in_buf[691]*(38)+in_buf[692]*(33)+in_buf[693]*(6)+in_buf[694]*(0)+in_buf[695]*(16)+in_buf[696]*(-16)+in_buf[697]*(-10)+in_buf[698]*(-11)+in_buf[699]*(-3)+in_buf[700]*(-3)+in_buf[701]*(0)+in_buf[702]*(-20)+in_buf[703]*(-25)+in_buf[704]*(-38)+in_buf[705]*(-7)+in_buf[706]*(14)+in_buf[707]*(17)+in_buf[708]*(17)+in_buf[709]*(20)+in_buf[710]*(16)+in_buf[711]*(-1)+in_buf[712]*(7)+in_buf[713]*(26)+in_buf[714]*(30)+in_buf[715]*(20)+in_buf[716]*(17)+in_buf[717]*(31)+in_buf[718]*(34)+in_buf[719]*(48)+in_buf[720]*(35)+in_buf[721]*(36)+in_buf[722]*(-4)+in_buf[723]*(1)+in_buf[724]*(-5)+in_buf[725]*(0)+in_buf[726]*(-11)+in_buf[727]*(1)+in_buf[728]*(-3)+in_buf[729]*(3)+in_buf[730]*(-2)+in_buf[731]*(4)+in_buf[732]*(26)+in_buf[733]*(39)+in_buf[734]*(38)+in_buf[735]*(26)+in_buf[736]*(22)+in_buf[737]*(23)+in_buf[738]*(19)+in_buf[739]*(9)+in_buf[740]*(19)+in_buf[741]*(27)+in_buf[742]*(50)+in_buf[743]*(34)+in_buf[744]*(33)+in_buf[745]*(52)+in_buf[746]*(44)+in_buf[747]*(0)+in_buf[748]*(24)+in_buf[749]*(43)+in_buf[750]*(18)+in_buf[751]*(25)+in_buf[752]*(21)+in_buf[753]*(-6)+in_buf[754]*(1)+in_buf[755]*(3)+in_buf[756]*(4)+in_buf[757]*(-1)+in_buf[758]*(3)+in_buf[759]*(2)+in_buf[760]*(-15)+in_buf[761]*(-34)+in_buf[762]*(6)+in_buf[763]*(6)+in_buf[764]*(8)+in_buf[765]*(0)+in_buf[766]*(1)+in_buf[767]*(24)+in_buf[768]*(23)+in_buf[769]*(0)+in_buf[770]*(37)+in_buf[771]*(34)+in_buf[772]*(-1)+in_buf[773]*(-14)+in_buf[774]*(3)+in_buf[775]*(23)+in_buf[776]*(8)+in_buf[777]*(-10)+in_buf[778]*(3)+in_buf[779]*(9)+in_buf[780]*(4)+in_buf[781]*(1)+in_buf[782]*(3)+in_buf[783]*(2);
assign in_buf_weight05=in_buf[0]*(-3)+in_buf[1]*(0)+in_buf[2]*(0)+in_buf[3]*(-1)+in_buf[4]*(0)+in_buf[5]*(4)+in_buf[6]*(4)+in_buf[7]*(0)+in_buf[8]*(2)+in_buf[9]*(0)+in_buf[10]*(-1)+in_buf[11]*(-3)+in_buf[12]*(-2)+in_buf[13]*(3)+in_buf[14]*(4)+in_buf[15]*(-2)+in_buf[16]*(1)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(-1)+in_buf[20]*(-1)+in_buf[21]*(4)+in_buf[22]*(3)+in_buf[23]*(-2)+in_buf[24]*(0)+in_buf[25]*(2)+in_buf[26]*(3)+in_buf[27]*(-3)+in_buf[28]*(-3)+in_buf[29]*(-3)+in_buf[30]*(0)+in_buf[31]*(0)+in_buf[32]*(4)+in_buf[33]*(0)+in_buf[34]*(-1)+in_buf[35]*(1)+in_buf[36]*(0)+in_buf[37]*(4)+in_buf[38]*(1)+in_buf[39]*(25)+in_buf[40]*(24)+in_buf[41]*(19)+in_buf[42]*(9)+in_buf[43]*(34)+in_buf[44]*(28)+in_buf[45]*(28)+in_buf[46]*(17)+in_buf[47]*(15)+in_buf[48]*(22)+in_buf[49]*(28)+in_buf[50]*(10)+in_buf[51]*(0)+in_buf[52]*(0)+in_buf[53]*(3)+in_buf[54]*(0)+in_buf[55]*(1)+in_buf[56]*(3)+in_buf[57]*(-1)+in_buf[58]*(10)+in_buf[59]*(10)+in_buf[60]*(18)+in_buf[61]*(5)+in_buf[62]*(14)+in_buf[63]*(25)+in_buf[64]*(-1)+in_buf[65]*(-11)+in_buf[66]*(-15)+in_buf[67]*(-1)+in_buf[68]*(-3)+in_buf[69]*(-37)+in_buf[70]*(-38)+in_buf[71]*(-9)+in_buf[72]*(7)+in_buf[73]*(8)+in_buf[74]*(15)+in_buf[75]*(4)+in_buf[76]*(1)+in_buf[77]*(7)+in_buf[78]*(34)+in_buf[79]*(9)+in_buf[80]*(-9)+in_buf[81]*(-5)+in_buf[82]*(-2)+in_buf[83]*(3)+in_buf[84]*(-3)+in_buf[85]*(-3)+in_buf[86]*(-2)+in_buf[87]*(7)+in_buf[88]*(23)+in_buf[89]*(11)+in_buf[90]*(12)+in_buf[91]*(7)+in_buf[92]*(-4)+in_buf[93]*(-29)+in_buf[94]*(-19)+in_buf[95]*(-32)+in_buf[96]*(-22)+in_buf[97]*(-24)+in_buf[98]*(-5)+in_buf[99]*(7)+in_buf[100]*(-1)+in_buf[101]*(27)+in_buf[102]*(37)+in_buf[103]*(0)+in_buf[104]*(14)+in_buf[105]*(18)+in_buf[106]*(16)+in_buf[107]*(58)+in_buf[108]*(19)+in_buf[109]*(-19)+in_buf[110]*(-18)+in_buf[111]*(-2)+in_buf[112]*(2)+in_buf[113]*(0)+in_buf[114]*(13)+in_buf[115]*(22)+in_buf[116]*(6)+in_buf[117]*(-10)+in_buf[118]*(-19)+in_buf[119]*(-15)+in_buf[120]*(-20)+in_buf[121]*(-8)+in_buf[122]*(-9)+in_buf[123]*(-7)+in_buf[124]*(-9)+in_buf[125]*(-16)+in_buf[126]*(-7)+in_buf[127]*(15)+in_buf[128]*(6)+in_buf[129]*(6)+in_buf[130]*(4)+in_buf[131]*(2)+in_buf[132]*(5)+in_buf[133]*(15)+in_buf[134]*(13)+in_buf[135]*(7)+in_buf[136]*(-17)+in_buf[137]*(9)+in_buf[138]*(31)+in_buf[139]*(18)+in_buf[140]*(0)+in_buf[141]*(4)+in_buf[142]*(43)+in_buf[143]*(6)+in_buf[144]*(-16)+in_buf[145]*(-9)+in_buf[146]*(-3)+in_buf[147]*(-1)+in_buf[148]*(-6)+in_buf[149]*(0)+in_buf[150]*(8)+in_buf[151]*(-5)+in_buf[152]*(-16)+in_buf[153]*(0)+in_buf[154]*(0)+in_buf[155]*(-6)+in_buf[156]*(-6)+in_buf[157]*(5)+in_buf[158]*(11)+in_buf[159]*(13)+in_buf[160]*(32)+in_buf[161]*(22)+in_buf[162]*(8)+in_buf[163]*(-22)+in_buf[164]*(-10)+in_buf[165]*(1)+in_buf[166]*(40)+in_buf[167]*(19)+in_buf[168]*(2)+in_buf[169]*(21)+in_buf[170]*(1)+in_buf[171]*(-9)+in_buf[172]*(-15)+in_buf[173]*(0)+in_buf[174]*(-5)+in_buf[175]*(10)+in_buf[176]*(24)+in_buf[177]*(4)+in_buf[178]*(-2)+in_buf[179]*(-15)+in_buf[180]*(-15)+in_buf[181]*(-7)+in_buf[182]*(-15)+in_buf[183]*(-13)+in_buf[184]*(-9)+in_buf[185]*(10)+in_buf[186]*(14)+in_buf[187]*(16)+in_buf[188]*(23)+in_buf[189]*(16)+in_buf[190]*(9)+in_buf[191]*(2)+in_buf[192]*(18)+in_buf[193]*(24)+in_buf[194]*(16)+in_buf[195]*(-5)+in_buf[196]*(-1)+in_buf[197]*(16)+in_buf[198]*(-5)+in_buf[199]*(-20)+in_buf[200]*(-29)+in_buf[201]*(5)+in_buf[202]*(-16)+in_buf[203]*(-3)+in_buf[204]*(5)+in_buf[205]*(-7)+in_buf[206]*(-15)+in_buf[207]*(-8)+in_buf[208]*(-13)+in_buf[209]*(-12)+in_buf[210]*(-17)+in_buf[211]*(14)+in_buf[212]*(10)+in_buf[213]*(16)+in_buf[214]*(32)+in_buf[215]*(24)+in_buf[216]*(24)+in_buf[217]*(13)+in_buf[218]*(19)+in_buf[219]*(22)+in_buf[220]*(9)+in_buf[221]*(28)+in_buf[222]*(-3)+in_buf[223]*(-9)+in_buf[224]*(1)+in_buf[225]*(6)+in_buf[226]*(-26)+in_buf[227]*(-6)+in_buf[228]*(-10)+in_buf[229]*(-3)+in_buf[230]*(12)+in_buf[231]*(3)+in_buf[232]*(-8)+in_buf[233]*(-10)+in_buf[234]*(-9)+in_buf[235]*(-7)+in_buf[236]*(5)+in_buf[237]*(0)+in_buf[238]*(-7)+in_buf[239]*(3)+in_buf[240]*(23)+in_buf[241]*(9)+in_buf[242]*(14)+in_buf[243]*(17)+in_buf[244]*(25)+in_buf[245]*(24)+in_buf[246]*(23)+in_buf[247]*(18)+in_buf[248]*(22)+in_buf[249]*(10)+in_buf[250]*(-9)+in_buf[251]*(7)+in_buf[252]*(-11)+in_buf[253]*(-5)+in_buf[254]*(-38)+in_buf[255]*(-16)+in_buf[256]*(-25)+in_buf[257]*(-13)+in_buf[258]*(10)+in_buf[259]*(-4)+in_buf[260]*(-10)+in_buf[261]*(4)+in_buf[262]*(12)+in_buf[263]*(4)+in_buf[264]*(-3)+in_buf[265]*(-1)+in_buf[266]*(-13)+in_buf[267]*(-11)+in_buf[268]*(2)+in_buf[269]*(-8)+in_buf[270]*(-11)+in_buf[271]*(0)+in_buf[272]*(10)+in_buf[273]*(14)+in_buf[274]*(21)+in_buf[275]*(31)+in_buf[276]*(35)+in_buf[277]*(36)+in_buf[278]*(-9)+in_buf[279]*(-18)+in_buf[280]*(-9)+in_buf[281]*(1)+in_buf[282]*(26)+in_buf[283]*(-12)+in_buf[284]*(-28)+in_buf[285]*(-18)+in_buf[286]*(-13)+in_buf[287]*(-10)+in_buf[288]*(-11)+in_buf[289]*(2)+in_buf[290]*(9)+in_buf[291]*(8)+in_buf[292]*(5)+in_buf[293]*(0)+in_buf[294]*(8)+in_buf[295]*(17)+in_buf[296]*(5)+in_buf[297]*(-11)+in_buf[298]*(0)+in_buf[299]*(-15)+in_buf[300]*(7)+in_buf[301]*(-3)+in_buf[302]*(21)+in_buf[303]*(42)+in_buf[304]*(39)+in_buf[305]*(14)+in_buf[306]*(12)+in_buf[307]*(-20)+in_buf[308]*(-7)+in_buf[309]*(-29)+in_buf[310]*(23)+in_buf[311]*(-3)+in_buf[312]*(-23)+in_buf[313]*(-11)+in_buf[314]*(0)+in_buf[315]*(0)+in_buf[316]*(-6)+in_buf[317]*(4)+in_buf[318]*(-1)+in_buf[319]*(6)+in_buf[320]*(4)+in_buf[321]*(34)+in_buf[322]*(42)+in_buf[323]*(34)+in_buf[324]*(4)+in_buf[325]*(4)+in_buf[326]*(3)+in_buf[327]*(-18)+in_buf[328]*(-16)+in_buf[329]*(-3)+in_buf[330]*(-8)+in_buf[331]*(17)+in_buf[332]*(24)+in_buf[333]*(20)+in_buf[334]*(54)+in_buf[335]*(-19)+in_buf[336]*(-2)+in_buf[337]*(-10)+in_buf[338]*(2)+in_buf[339]*(-1)+in_buf[340]*(-15)+in_buf[341]*(-1)+in_buf[342]*(0)+in_buf[343]*(-4)+in_buf[344]*(-12)+in_buf[345]*(8)+in_buf[346]*(2)+in_buf[347]*(12)+in_buf[348]*(5)+in_buf[349]*(35)+in_buf[350]*(53)+in_buf[351]*(33)+in_buf[352]*(0)+in_buf[353]*(11)+in_buf[354]*(1)+in_buf[355]*(-22)+in_buf[356]*(-15)+in_buf[357]*(-17)+in_buf[358]*(-16)+in_buf[359]*(-15)+in_buf[360]*(-24)+in_buf[361]*(-18)+in_buf[362]*(10)+in_buf[363]*(-32)+in_buf[364]*(15)+in_buf[365]*(-4)+in_buf[366]*(-27)+in_buf[367]*(-18)+in_buf[368]*(-17)+in_buf[369]*(8)+in_buf[370]*(3)+in_buf[371]*(-13)+in_buf[372]*(-3)+in_buf[373]*(6)+in_buf[374]*(0)+in_buf[375]*(9)+in_buf[376]*(19)+in_buf[377]*(20)+in_buf[378]*(27)+in_buf[379]*(7)+in_buf[380]*(-13)+in_buf[381]*(-11)+in_buf[382]*(-26)+in_buf[383]*(-22)+in_buf[384]*(-28)+in_buf[385]*(-16)+in_buf[386]*(-20)+in_buf[387]*(0)+in_buf[388]*(-30)+in_buf[389]*(-22)+in_buf[390]*(-15)+in_buf[391]*(-10)+in_buf[392]*(14)+in_buf[393]*(-7)+in_buf[394]*(-25)+in_buf[395]*(-30)+in_buf[396]*(0)+in_buf[397]*(8)+in_buf[398]*(0)+in_buf[399]*(-17)+in_buf[400]*(4)+in_buf[401]*(7)+in_buf[402]*(8)+in_buf[403]*(13)+in_buf[404]*(14)+in_buf[405]*(17)+in_buf[406]*(12)+in_buf[407]*(-8)+in_buf[408]*(-18)+in_buf[409]*(-9)+in_buf[410]*(-16)+in_buf[411]*(-26)+in_buf[412]*(-9)+in_buf[413]*(0)+in_buf[414]*(-19)+in_buf[415]*(-4)+in_buf[416]*(2)+in_buf[417]*(-6)+in_buf[418]*(-37)+in_buf[419]*(-12)+in_buf[420]*(7)+in_buf[421]*(10)+in_buf[422]*(-21)+in_buf[423]*(-53)+in_buf[424]*(4)+in_buf[425]*(14)+in_buf[426]*(19)+in_buf[427]*(11)+in_buf[428]*(21)+in_buf[429]*(12)+in_buf[430]*(5)+in_buf[431]*(11)+in_buf[432]*(21)+in_buf[433]*(1)+in_buf[434]*(-8)+in_buf[435]*(-33)+in_buf[436]*(-8)+in_buf[437]*(-2)+in_buf[438]*(5)+in_buf[439]*(-13)+in_buf[440]*(-9)+in_buf[441]*(-19)+in_buf[442]*(-23)+in_buf[443]*(3)+in_buf[444]*(30)+in_buf[445]*(-13)+in_buf[446]*(-36)+in_buf[447]*(-14)+in_buf[448]*(-5)+in_buf[449]*(6)+in_buf[450]*(5)+in_buf[451]*(-27)+in_buf[452]*(-1)+in_buf[453]*(11)+in_buf[454]*(13)+in_buf[455]*(-2)+in_buf[456]*(17)+in_buf[457]*(20)+in_buf[458]*(18)+in_buf[459]*(19)+in_buf[460]*(2)+in_buf[461]*(-17)+in_buf[462]*(-31)+in_buf[463]*(-30)+in_buf[464]*(-8)+in_buf[465]*(-4)+in_buf[466]*(1)+in_buf[467]*(-5)+in_buf[468]*(-13)+in_buf[469]*(-36)+in_buf[470]*(-20)+in_buf[471]*(-21)+in_buf[472]*(22)+in_buf[473]*(-26)+in_buf[474]*(-55)+in_buf[475]*(-17)+in_buf[476]*(2)+in_buf[477]*(11)+in_buf[478]*(-24)+in_buf[479]*(2)+in_buf[480]*(0)+in_buf[481]*(6)+in_buf[482]*(9)+in_buf[483]*(3)+in_buf[484]*(5)+in_buf[485]*(7)+in_buf[486]*(8)+in_buf[487]*(-4)+in_buf[488]*(-22)+in_buf[489]*(-37)+in_buf[490]*(-30)+in_buf[491]*(-9)+in_buf[492]*(5)+in_buf[493]*(20)+in_buf[494]*(8)+in_buf[495]*(20)+in_buf[496]*(-3)+in_buf[497]*(-26)+in_buf[498]*(-33)+in_buf[499]*(-6)+in_buf[500]*(-5)+in_buf[501]*(-44)+in_buf[502]*(-45)+in_buf[503]*(13)+in_buf[504]*(35)+in_buf[505]*(13)+in_buf[506]*(-6)+in_buf[507]*(-10)+in_buf[508]*(-6)+in_buf[509]*(11)+in_buf[510]*(5)+in_buf[511]*(4)+in_buf[512]*(11)+in_buf[513]*(12)+in_buf[514]*(9)+in_buf[515]*(-9)+in_buf[516]*(-28)+in_buf[517]*(-28)+in_buf[518]*(-22)+in_buf[519]*(0)+in_buf[520]*(-1)+in_buf[521]*(18)+in_buf[522]*(15)+in_buf[523]*(2)+in_buf[524]*(0)+in_buf[525]*(-10)+in_buf[526]*(-41)+in_buf[527]*(-29)+in_buf[528]*(-21)+in_buf[529]*(-19)+in_buf[530]*(-39)+in_buf[531]*(-26)+in_buf[532]*(1)+in_buf[533]*(43)+in_buf[534]*(8)+in_buf[535]*(-25)+in_buf[536]*(-11)+in_buf[537]*(7)+in_buf[538]*(20)+in_buf[539]*(-2)+in_buf[540]*(14)+in_buf[541]*(16)+in_buf[542]*(12)+in_buf[543]*(-9)+in_buf[544]*(-3)+in_buf[545]*(-24)+in_buf[546]*(-29)+in_buf[547]*(-11)+in_buf[548]*(-1)+in_buf[549]*(16)+in_buf[550]*(21)+in_buf[551]*(0)+in_buf[552]*(0)+in_buf[553]*(-24)+in_buf[554]*(-31)+in_buf[555]*(-8)+in_buf[556]*(16)+in_buf[557]*(-1)+in_buf[558]*(-27)+in_buf[559]*(-25)+in_buf[560]*(4)+in_buf[561]*(29)+in_buf[562]*(-23)+in_buf[563]*(-32)+in_buf[564]*(-1)+in_buf[565]*(9)+in_buf[566]*(0)+in_buf[567]*(0)+in_buf[568]*(19)+in_buf[569]*(18)+in_buf[570]*(21)+in_buf[571]*(7)+in_buf[572]*(10)+in_buf[573]*(0)+in_buf[574]*(-19)+in_buf[575]*(-4)+in_buf[576]*(-3)+in_buf[577]*(15)+in_buf[578]*(5)+in_buf[579]*(-7)+in_buf[580]*(0)+in_buf[581]*(-15)+in_buf[582]*(-16)+in_buf[583]*(-22)+in_buf[584]*(6)+in_buf[585]*(-5)+in_buf[586]*(-12)+in_buf[587]*(10)+in_buf[588]*(-15)+in_buf[589]*(8)+in_buf[590]*(-24)+in_buf[591]*(-23)+in_buf[592]*(-8)+in_buf[593]*(-7)+in_buf[594]*(4)+in_buf[595]*(6)+in_buf[596]*(5)+in_buf[597]*(12)+in_buf[598]*(7)+in_buf[599]*(18)+in_buf[600]*(9)+in_buf[601]*(0)+in_buf[602]*(-10)+in_buf[603]*(2)+in_buf[604]*(5)+in_buf[605]*(13)+in_buf[606]*(0)+in_buf[607]*(0)+in_buf[608]*(-1)+in_buf[609]*(-12)+in_buf[610]*(-35)+in_buf[611]*(-25)+in_buf[612]*(0)+in_buf[613]*(-3)+in_buf[614]*(12)+in_buf[615]*(0)+in_buf[616]*(-9)+in_buf[617]*(2)+in_buf[618]*(-13)+in_buf[619]*(2)+in_buf[620]*(-7)+in_buf[621]*(-2)+in_buf[622]*(2)+in_buf[623]*(4)+in_buf[624]*(-8)+in_buf[625]*(10)+in_buf[626]*(13)+in_buf[627]*(29)+in_buf[628]*(19)+in_buf[629]*(10)+in_buf[630]*(1)+in_buf[631]*(6)+in_buf[632]*(6)+in_buf[633]*(-9)+in_buf[634]*(-24)+in_buf[635]*(-14)+in_buf[636]*(-20)+in_buf[637]*(-30)+in_buf[638]*(-25)+in_buf[639]*(-24)+in_buf[640]*(-22)+in_buf[641]*(-3)+in_buf[642]*(-5)+in_buf[643]*(-2)+in_buf[644]*(-2)+in_buf[645]*(-1)+in_buf[646]*(28)+in_buf[647]*(27)+in_buf[648]*(13)+in_buf[649]*(-4)+in_buf[650]*(-10)+in_buf[651]*(0)+in_buf[652]*(1)+in_buf[653]*(-1)+in_buf[654]*(1)+in_buf[655]*(25)+in_buf[656]*(25)+in_buf[657]*(26)+in_buf[658]*(2)+in_buf[659]*(15)+in_buf[660]*(-6)+in_buf[661]*(-21)+in_buf[662]*(-43)+in_buf[663]*(-41)+in_buf[664]*(-26)+in_buf[665]*(-18)+in_buf[666]*(-19)+in_buf[667]*(-20)+in_buf[668]*(-17)+in_buf[669]*(-9)+in_buf[670]*(-20)+in_buf[671]*(-2)+in_buf[672]*(-3)+in_buf[673]*(1)+in_buf[674]*(11)+in_buf[675]*(30)+in_buf[676]*(10)+in_buf[677]*(10)+in_buf[678]*(-9)+in_buf[679]*(-6)+in_buf[680]*(16)+in_buf[681]*(19)+in_buf[682]*(20)+in_buf[683]*(13)+in_buf[684]*(38)+in_buf[685]*(17)+in_buf[686]*(3)+in_buf[687]*(17)+in_buf[688]*(12)+in_buf[689]*(-17)+in_buf[690]*(-35)+in_buf[691]*(-37)+in_buf[692]*(-1)+in_buf[693]*(-22)+in_buf[694]*(-25)+in_buf[695]*(-27)+in_buf[696]*(-8)+in_buf[697]*(-30)+in_buf[698]*(-9)+in_buf[699]*(-1)+in_buf[700]*(-1)+in_buf[701]*(1)+in_buf[702]*(8)+in_buf[703]*(10)+in_buf[704]*(-29)+in_buf[705]*(0)+in_buf[706]*(25)+in_buf[707]*(33)+in_buf[708]*(16)+in_buf[709]*(20)+in_buf[710]*(16)+in_buf[711]*(12)+in_buf[712]*(9)+in_buf[713]*(3)+in_buf[714]*(-2)+in_buf[715]*(11)+in_buf[716]*(16)+in_buf[717]*(0)+in_buf[718]*(-10)+in_buf[719]*(13)+in_buf[720]*(4)+in_buf[721]*(2)+in_buf[722]*(9)+in_buf[723]*(-9)+in_buf[724]*(-6)+in_buf[725]*(-5)+in_buf[726]*(-3)+in_buf[727]*(0)+in_buf[728]*(2)+in_buf[729]*(3)+in_buf[730]*(3)+in_buf[731]*(4)+in_buf[732]*(32)+in_buf[733]*(34)+in_buf[734]*(7)+in_buf[735]*(-1)+in_buf[736]*(21)+in_buf[737]*(12)+in_buf[738]*(27)+in_buf[739]*(36)+in_buf[740]*(29)+in_buf[741]*(15)+in_buf[742]*(18)+in_buf[743]*(0)+in_buf[744]*(21)+in_buf[745]*(18)+in_buf[746]*(6)+in_buf[747]*(11)+in_buf[748]*(24)+in_buf[749]*(22)+in_buf[750]*(9)+in_buf[751]*(2)+in_buf[752]*(4)+in_buf[753]*(3)+in_buf[754]*(-2)+in_buf[755]*(2)+in_buf[756]*(4)+in_buf[757]*(-2)+in_buf[758]*(-1)+in_buf[759]*(4)+in_buf[760]*(-20)+in_buf[761]*(-18)+in_buf[762]*(-1)+in_buf[763]*(6)+in_buf[764]*(3)+in_buf[765]*(-16)+in_buf[766]*(15)+in_buf[767]*(8)+in_buf[768]*(6)+in_buf[769]*(-11)+in_buf[770]*(27)+in_buf[771]*(21)+in_buf[772]*(22)+in_buf[773]*(-1)+in_buf[774]*(6)+in_buf[775]*(0)+in_buf[776]*(0)+in_buf[777]*(-4)+in_buf[778]*(-7)+in_buf[779]*(-3)+in_buf[780]*(3)+in_buf[781]*(1)+in_buf[782]*(0)+in_buf[783]*(-1);
assign in_buf_weight06=in_buf[0]*(4)+in_buf[1]*(-1)+in_buf[2]*(4)+in_buf[3]*(1)+in_buf[4]*(2)+in_buf[5]*(3)+in_buf[6]*(-1)+in_buf[7]*(4)+in_buf[8]*(2)+in_buf[9]*(-3)+in_buf[10]*(-1)+in_buf[11]*(3)+in_buf[12]*(0)+in_buf[13]*(2)+in_buf[14]*(4)+in_buf[15]*(4)+in_buf[16]*(0)+in_buf[17]*(-2)+in_buf[18]*(1)+in_buf[19]*(-1)+in_buf[20]*(1)+in_buf[21]*(1)+in_buf[22]*(0)+in_buf[23]*(0)+in_buf[24]*(4)+in_buf[25]*(-3)+in_buf[26]*(4)+in_buf[27]*(0)+in_buf[28]*(0)+in_buf[29]*(-1)+in_buf[30]*(5)+in_buf[31]*(-1)+in_buf[32]*(2)+in_buf[33]*(0)+in_buf[34]*(-1)+in_buf[35]*(-3)+in_buf[36]*(-1)+in_buf[37]*(1)+in_buf[38]*(2)+in_buf[39]*(1)+in_buf[40]*(4)+in_buf[41]*(-3)+in_buf[42]*(1)+in_buf[43]*(3)+in_buf[44]*(4)+in_buf[45]*(-2)+in_buf[46]*(-3)+in_buf[47]*(0)+in_buf[48]*(-3)+in_buf[49]*(0)+in_buf[50]*(0)+in_buf[51]*(-1)+in_buf[52]*(1)+in_buf[53]*(-1)+in_buf[54]*(2)+in_buf[55]*(1)+in_buf[56]*(-3)+in_buf[57]*(-1)+in_buf[58]*(-2)+in_buf[59]*(4)+in_buf[60]*(4)+in_buf[61]*(-1)+in_buf[62]*(-1)+in_buf[63]*(3)+in_buf[64]*(-2)+in_buf[65]*(1)+in_buf[66]*(1)+in_buf[67]*(1)+in_buf[68]*(-3)+in_buf[69]*(-3)+in_buf[70]*(2)+in_buf[71]*(-1)+in_buf[72]*(-3)+in_buf[73]*(-1)+in_buf[74]*(-2)+in_buf[75]*(3)+in_buf[76]*(1)+in_buf[77]*(3)+in_buf[78]*(-2)+in_buf[79]*(0)+in_buf[80]*(0)+in_buf[81]*(4)+in_buf[82]*(4)+in_buf[83]*(1)+in_buf[84]*(0)+in_buf[85]*(-3)+in_buf[86]*(-1)+in_buf[87]*(-3)+in_buf[88]*(4)+in_buf[89]*(-3)+in_buf[90]*(2)+in_buf[91]*(4)+in_buf[92]*(1)+in_buf[93]*(-1)+in_buf[94]*(-5)+in_buf[95]*(0)+in_buf[96]*(1)+in_buf[97]*(0)+in_buf[98]*(-2)+in_buf[99]*(0)+in_buf[100]*(-1)+in_buf[101]*(4)+in_buf[102]*(-2)+in_buf[103]*(3)+in_buf[104]*(-3)+in_buf[105]*(0)+in_buf[106]*(-1)+in_buf[107]*(-3)+in_buf[108]*(2)+in_buf[109]*(2)+in_buf[110]*(3)+in_buf[111]*(-1)+in_buf[112]*(-1)+in_buf[113]*(2)+in_buf[114]*(-2)+in_buf[115]*(0)+in_buf[116]*(-3)+in_buf[117]*(-3)+in_buf[118]*(-3)+in_buf[119]*(0)+in_buf[120]*(-5)+in_buf[121]*(-1)+in_buf[122]*(-2)+in_buf[123]*(2)+in_buf[124]*(-3)+in_buf[125]*(0)+in_buf[126]*(-1)+in_buf[127]*(1)+in_buf[128]*(-3)+in_buf[129]*(1)+in_buf[130]*(-3)+in_buf[131]*(-4)+in_buf[132]*(2)+in_buf[133]*(-3)+in_buf[134]*(1)+in_buf[135]*(3)+in_buf[136]*(0)+in_buf[137]*(2)+in_buf[138]*(4)+in_buf[139]*(0)+in_buf[140]*(2)+in_buf[141]*(2)+in_buf[142]*(1)+in_buf[143]*(-3)+in_buf[144]*(3)+in_buf[145]*(0)+in_buf[146]*(-3)+in_buf[147]*(0)+in_buf[148]*(0)+in_buf[149]*(3)+in_buf[150]*(-3)+in_buf[151]*(0)+in_buf[152]*(-2)+in_buf[153]*(-3)+in_buf[154]*(0)+in_buf[155]*(-2)+in_buf[156]*(-4)+in_buf[157]*(0)+in_buf[158]*(-3)+in_buf[159]*(-2)+in_buf[160]*(1)+in_buf[161]*(0)+in_buf[162]*(4)+in_buf[163]*(-1)+in_buf[164]*(1)+in_buf[165]*(1)+in_buf[166]*(0)+in_buf[167]*(0)+in_buf[168]*(0)+in_buf[169]*(4)+in_buf[170]*(-2)+in_buf[171]*(0)+in_buf[172]*(2)+in_buf[173]*(-1)+in_buf[174]*(-3)+in_buf[175]*(2)+in_buf[176]*(0)+in_buf[177]*(-1)+in_buf[178]*(0)+in_buf[179]*(-3)+in_buf[180]*(-3)+in_buf[181]*(-2)+in_buf[182]*(3)+in_buf[183]*(-4)+in_buf[184]*(0)+in_buf[185]*(-1)+in_buf[186]*(-1)+in_buf[187]*(-2)+in_buf[188]*(3)+in_buf[189]*(-2)+in_buf[190]*(-3)+in_buf[191]*(3)+in_buf[192]*(0)+in_buf[193]*(-2)+in_buf[194]*(0)+in_buf[195]*(4)+in_buf[196]*(0)+in_buf[197]*(1)+in_buf[198]*(2)+in_buf[199]*(3)+in_buf[200]*(4)+in_buf[201]*(3)+in_buf[202]*(1)+in_buf[203]*(1)+in_buf[204]*(0)+in_buf[205]*(-1)+in_buf[206]*(0)+in_buf[207]*(-2)+in_buf[208]*(-2)+in_buf[209]*(-3)+in_buf[210]*(3)+in_buf[211]*(-2)+in_buf[212]*(-4)+in_buf[213]*(0)+in_buf[214]*(-3)+in_buf[215]*(2)+in_buf[216]*(1)+in_buf[217]*(0)+in_buf[218]*(-2)+in_buf[219]*(0)+in_buf[220]*(0)+in_buf[221]*(2)+in_buf[222]*(-3)+in_buf[223]*(3)+in_buf[224]*(0)+in_buf[225]*(-3)+in_buf[226]*(4)+in_buf[227]*(-1)+in_buf[228]*(-2)+in_buf[229]*(2)+in_buf[230]*(-2)+in_buf[231]*(2)+in_buf[232]*(0)+in_buf[233]*(-3)+in_buf[234]*(-1)+in_buf[235]*(0)+in_buf[236]*(-3)+in_buf[237]*(-3)+in_buf[238]*(2)+in_buf[239]*(3)+in_buf[240]*(-4)+in_buf[241]*(0)+in_buf[242]*(0)+in_buf[243]*(-3)+in_buf[244]*(1)+in_buf[245]*(3)+in_buf[246]*(-3)+in_buf[247]*(3)+in_buf[248]*(1)+in_buf[249]*(0)+in_buf[250]*(-2)+in_buf[251]*(0)+in_buf[252]*(3)+in_buf[253]*(0)+in_buf[254]*(2)+in_buf[255]*(2)+in_buf[256]*(-2)+in_buf[257]*(-3)+in_buf[258]*(-1)+in_buf[259]*(2)+in_buf[260]*(-1)+in_buf[261]*(-1)+in_buf[262]*(0)+in_buf[263]*(2)+in_buf[264]*(1)+in_buf[265]*(0)+in_buf[266]*(-1)+in_buf[267]*(-3)+in_buf[268]*(2)+in_buf[269]*(-3)+in_buf[270]*(3)+in_buf[271]*(-4)+in_buf[272]*(1)+in_buf[273]*(0)+in_buf[274]*(0)+in_buf[275]*(0)+in_buf[276]*(1)+in_buf[277]*(4)+in_buf[278]*(0)+in_buf[279]*(4)+in_buf[280]*(0)+in_buf[281]*(-2)+in_buf[282]*(3)+in_buf[283]*(3)+in_buf[284]*(-2)+in_buf[285]*(-4)+in_buf[286]*(-4)+in_buf[287]*(-2)+in_buf[288]*(-2)+in_buf[289]*(2)+in_buf[290]*(0)+in_buf[291]*(-4)+in_buf[292]*(2)+in_buf[293]*(1)+in_buf[294]*(3)+in_buf[295]*(0)+in_buf[296]*(3)+in_buf[297]*(-4)+in_buf[298]*(0)+in_buf[299]*(-3)+in_buf[300]*(1)+in_buf[301]*(-1)+in_buf[302]*(0)+in_buf[303]*(-1)+in_buf[304]*(-4)+in_buf[305]*(-2)+in_buf[306]*(1)+in_buf[307]*(3)+in_buf[308]*(0)+in_buf[309]*(-2)+in_buf[310]*(-1)+in_buf[311]*(-1)+in_buf[312]*(-1)+in_buf[313]*(0)+in_buf[314]*(-3)+in_buf[315]*(4)+in_buf[316]*(2)+in_buf[317]*(-2)+in_buf[318]*(-4)+in_buf[319]*(1)+in_buf[320]*(-4)+in_buf[321]*(-4)+in_buf[322]*(-2)+in_buf[323]*(0)+in_buf[324]*(0)+in_buf[325]*(0)+in_buf[326]*(-1)+in_buf[327]*(4)+in_buf[328]*(0)+in_buf[329]*(0)+in_buf[330]*(3)+in_buf[331]*(-4)+in_buf[332]*(2)+in_buf[333]*(3)+in_buf[334]*(0)+in_buf[335]*(4)+in_buf[336]*(-3)+in_buf[337]*(3)+in_buf[338]*(0)+in_buf[339]*(-2)+in_buf[340]*(2)+in_buf[341]*(0)+in_buf[342]*(1)+in_buf[343]*(0)+in_buf[344]*(-1)+in_buf[345]*(-3)+in_buf[346]*(-1)+in_buf[347]*(-4)+in_buf[348]*(-2)+in_buf[349]*(3)+in_buf[350]*(2)+in_buf[351]*(-4)+in_buf[352]*(-3)+in_buf[353]*(2)+in_buf[354]*(2)+in_buf[355]*(3)+in_buf[356]*(3)+in_buf[357]*(-1)+in_buf[358]*(2)+in_buf[359]*(-1)+in_buf[360]*(-4)+in_buf[361]*(3)+in_buf[362]*(-3)+in_buf[363]*(1)+in_buf[364]*(0)+in_buf[365]*(2)+in_buf[366]*(1)+in_buf[367]*(3)+in_buf[368]*(0)+in_buf[369]*(-3)+in_buf[370]*(2)+in_buf[371]*(-1)+in_buf[372]*(-1)+in_buf[373]*(0)+in_buf[374]*(-4)+in_buf[375]*(-3)+in_buf[376]*(1)+in_buf[377]*(0)+in_buf[378]*(0)+in_buf[379]*(0)+in_buf[380]*(3)+in_buf[381]*(3)+in_buf[382]*(-3)+in_buf[383]*(-1)+in_buf[384]*(1)+in_buf[385]*(-3)+in_buf[386]*(0)+in_buf[387]*(-1)+in_buf[388]*(0)+in_buf[389]*(0)+in_buf[390]*(4)+in_buf[391]*(-1)+in_buf[392]*(0)+in_buf[393]*(0)+in_buf[394]*(3)+in_buf[395]*(1)+in_buf[396]*(-2)+in_buf[397]*(2)+in_buf[398]*(-3)+in_buf[399]*(0)+in_buf[400]*(2)+in_buf[401]*(-2)+in_buf[402]*(-4)+in_buf[403]*(0)+in_buf[404]*(2)+in_buf[405]*(-3)+in_buf[406]*(0)+in_buf[407]*(0)+in_buf[408]*(1)+in_buf[409]*(-1)+in_buf[410]*(-1)+in_buf[411]*(-1)+in_buf[412]*(-2)+in_buf[413]*(-2)+in_buf[414]*(1)+in_buf[415]*(2)+in_buf[416]*(-3)+in_buf[417]*(2)+in_buf[418]*(0)+in_buf[419]*(2)+in_buf[420]*(0)+in_buf[421]*(3)+in_buf[422]*(0)+in_buf[423]*(4)+in_buf[424]*(0)+in_buf[425]*(-2)+in_buf[426]*(1)+in_buf[427]*(3)+in_buf[428]*(-4)+in_buf[429]*(-2)+in_buf[430]*(0)+in_buf[431]*(-3)+in_buf[432]*(-1)+in_buf[433]*(-4)+in_buf[434]*(-3)+in_buf[435]*(-3)+in_buf[436]*(0)+in_buf[437]*(0)+in_buf[438]*(-1)+in_buf[439]*(3)+in_buf[440]*(3)+in_buf[441]*(0)+in_buf[442]*(-1)+in_buf[443]*(2)+in_buf[444]*(-2)+in_buf[445]*(-3)+in_buf[446]*(4)+in_buf[447]*(1)+in_buf[448]*(1)+in_buf[449]*(0)+in_buf[450]*(0)+in_buf[451]*(0)+in_buf[452]*(0)+in_buf[453]*(-1)+in_buf[454]*(-2)+in_buf[455]*(1)+in_buf[456]*(2)+in_buf[457]*(3)+in_buf[458]*(0)+in_buf[459]*(0)+in_buf[460]*(-4)+in_buf[461]*(1)+in_buf[462]*(2)+in_buf[463]*(-3)+in_buf[464]*(1)+in_buf[465]*(0)+in_buf[466]*(2)+in_buf[467]*(-3)+in_buf[468]*(-1)+in_buf[469]*(-2)+in_buf[470]*(-4)+in_buf[471]*(2)+in_buf[472]*(4)+in_buf[473]*(-3)+in_buf[474]*(1)+in_buf[475]*(-3)+in_buf[476]*(0)+in_buf[477]*(-2)+in_buf[478]*(-1)+in_buf[479]*(0)+in_buf[480]*(3)+in_buf[481]*(1)+in_buf[482]*(-3)+in_buf[483]*(-3)+in_buf[484]*(1)+in_buf[485]*(0)+in_buf[486]*(-3)+in_buf[487]*(3)+in_buf[488]*(-4)+in_buf[489]*(-2)+in_buf[490]*(1)+in_buf[491]*(0)+in_buf[492]*(-2)+in_buf[493]*(-3)+in_buf[494]*(-2)+in_buf[495]*(0)+in_buf[496]*(-3)+in_buf[497]*(2)+in_buf[498]*(-4)+in_buf[499]*(-2)+in_buf[500]*(0)+in_buf[501]*(4)+in_buf[502]*(-4)+in_buf[503]*(2)+in_buf[504]*(-1)+in_buf[505]*(2)+in_buf[506]*(-2)+in_buf[507]*(-2)+in_buf[508]*(1)+in_buf[509]*(1)+in_buf[510]*(-1)+in_buf[511]*(3)+in_buf[512]*(3)+in_buf[513]*(-4)+in_buf[514]*(-1)+in_buf[515]*(-2)+in_buf[516]*(-3)+in_buf[517]*(-4)+in_buf[518]*(4)+in_buf[519]*(0)+in_buf[520]*(-4)+in_buf[521]*(0)+in_buf[522]*(0)+in_buf[523]*(3)+in_buf[524]*(-1)+in_buf[525]*(-1)+in_buf[526]*(-3)+in_buf[527]*(0)+in_buf[528]*(2)+in_buf[529]*(-3)+in_buf[530]*(2)+in_buf[531]*(0)+in_buf[532]*(-3)+in_buf[533]*(0)+in_buf[534]*(1)+in_buf[535]*(3)+in_buf[536]*(0)+in_buf[537]*(0)+in_buf[538]*(-2)+in_buf[539]*(2)+in_buf[540]*(-2)+in_buf[541]*(0)+in_buf[542]*(-4)+in_buf[543]*(3)+in_buf[544]*(1)+in_buf[545]*(0)+in_buf[546]*(2)+in_buf[547]*(3)+in_buf[548]*(-1)+in_buf[549]*(3)+in_buf[550]*(-3)+in_buf[551]*(3)+in_buf[552]*(0)+in_buf[553]*(2)+in_buf[554]*(-3)+in_buf[555]*(0)+in_buf[556]*(1)+in_buf[557]*(0)+in_buf[558]*(0)+in_buf[559]*(-3)+in_buf[560]*(3)+in_buf[561]*(-1)+in_buf[562]*(-2)+in_buf[563]*(-3)+in_buf[564]*(3)+in_buf[565]*(0)+in_buf[566]*(-5)+in_buf[567]*(-1)+in_buf[568]*(-1)+in_buf[569]*(2)+in_buf[570]*(0)+in_buf[571]*(-4)+in_buf[572]*(-5)+in_buf[573]*(0)+in_buf[574]*(-1)+in_buf[575]*(-2)+in_buf[576]*(-1)+in_buf[577]*(2)+in_buf[578]*(-2)+in_buf[579]*(2)+in_buf[580]*(2)+in_buf[581]*(-3)+in_buf[582]*(2)+in_buf[583]*(3)+in_buf[584]*(0)+in_buf[585]*(4)+in_buf[586]*(2)+in_buf[587]*(-2)+in_buf[588]*(0)+in_buf[589]*(0)+in_buf[590]*(0)+in_buf[591]*(1)+in_buf[592]*(5)+in_buf[593]*(1)+in_buf[594]*(-3)+in_buf[595]*(1)+in_buf[596]*(-4)+in_buf[597]*(2)+in_buf[598]*(2)+in_buf[599]*(1)+in_buf[600]*(0)+in_buf[601]*(3)+in_buf[602]*(0)+in_buf[603]*(2)+in_buf[604]*(2)+in_buf[605]*(-5)+in_buf[606]*(3)+in_buf[607]*(0)+in_buf[608]*(-1)+in_buf[609]*(2)+in_buf[610]*(2)+in_buf[611]*(1)+in_buf[612]*(-2)+in_buf[613]*(1)+in_buf[614]*(0)+in_buf[615]*(3)+in_buf[616]*(2)+in_buf[617]*(0)+in_buf[618]*(2)+in_buf[619]*(0)+in_buf[620]*(3)+in_buf[621]*(-1)+in_buf[622]*(3)+in_buf[623]*(-3)+in_buf[624]*(0)+in_buf[625]*(-2)+in_buf[626]*(-3)+in_buf[627]*(-4)+in_buf[628]*(3)+in_buf[629]*(3)+in_buf[630]*(2)+in_buf[631]*(-2)+in_buf[632]*(-4)+in_buf[633]*(0)+in_buf[634]*(-4)+in_buf[635]*(0)+in_buf[636]*(1)+in_buf[637]*(4)+in_buf[638]*(1)+in_buf[639]*(-2)+in_buf[640]*(0)+in_buf[641]*(0)+in_buf[642]*(0)+in_buf[643]*(0)+in_buf[644]*(1)+in_buf[645]*(4)+in_buf[646]*(4)+in_buf[647]*(-1)+in_buf[648]*(2)+in_buf[649]*(4)+in_buf[650]*(1)+in_buf[651]*(5)+in_buf[652]*(2)+in_buf[653]*(0)+in_buf[654]*(-1)+in_buf[655]*(3)+in_buf[656]*(-5)+in_buf[657]*(-2)+in_buf[658]*(-3)+in_buf[659]*(-2)+in_buf[660]*(4)+in_buf[661]*(-2)+in_buf[662]*(-1)+in_buf[663]*(5)+in_buf[664]*(0)+in_buf[665]*(1)+in_buf[666]*(3)+in_buf[667]*(0)+in_buf[668]*(1)+in_buf[669]*(0)+in_buf[670]*(-3)+in_buf[671]*(0)+in_buf[672]*(3)+in_buf[673]*(3)+in_buf[674]*(3)+in_buf[675]*(0)+in_buf[676]*(0)+in_buf[677]*(-2)+in_buf[678]*(0)+in_buf[679]*(-2)+in_buf[680]*(1)+in_buf[681]*(0)+in_buf[682]*(5)+in_buf[683]*(0)+in_buf[684]*(-2)+in_buf[685]*(-2)+in_buf[686]*(-1)+in_buf[687]*(-2)+in_buf[688]*(-1)+in_buf[689]*(-2)+in_buf[690]*(3)+in_buf[691]*(3)+in_buf[692]*(1)+in_buf[693]*(0)+in_buf[694]*(-1)+in_buf[695]*(-3)+in_buf[696]*(3)+in_buf[697]*(3)+in_buf[698]*(0)+in_buf[699]*(-2)+in_buf[700]*(-1)+in_buf[701]*(-3)+in_buf[702]*(1)+in_buf[703]*(2)+in_buf[704]*(-2)+in_buf[705]*(4)+in_buf[706]*(-3)+in_buf[707]*(4)+in_buf[708]*(2)+in_buf[709]*(3)+in_buf[710]*(-1)+in_buf[711]*(4)+in_buf[712]*(-1)+in_buf[713]*(0)+in_buf[714]*(0)+in_buf[715]*(-2)+in_buf[716]*(-2)+in_buf[717]*(5)+in_buf[718]*(0)+in_buf[719]*(1)+in_buf[720]*(-2)+in_buf[721]*(-1)+in_buf[722]*(2)+in_buf[723]*(3)+in_buf[724]*(2)+in_buf[725]*(1)+in_buf[726]*(-4)+in_buf[727]*(-1)+in_buf[728]*(2)+in_buf[729]*(-3)+in_buf[730]*(2)+in_buf[731]*(-1)+in_buf[732]*(-1)+in_buf[733]*(0)+in_buf[734]*(3)+in_buf[735]*(0)+in_buf[736]*(-1)+in_buf[737]*(0)+in_buf[738]*(3)+in_buf[739]*(1)+in_buf[740]*(2)+in_buf[741]*(1)+in_buf[742]*(1)+in_buf[743]*(1)+in_buf[744]*(-3)+in_buf[745]*(4)+in_buf[746]*(0)+in_buf[747]*(2)+in_buf[748]*(1)+in_buf[749]*(-2)+in_buf[750]*(1)+in_buf[751]*(4)+in_buf[752]*(-2)+in_buf[753]*(-1)+in_buf[754]*(2)+in_buf[755]*(-3)+in_buf[756]*(3)+in_buf[757]*(0)+in_buf[758]*(1)+in_buf[759]*(2)+in_buf[760]*(4)+in_buf[761]*(0)+in_buf[762]*(2)+in_buf[763]*(-2)+in_buf[764]*(0)+in_buf[765]*(1)+in_buf[766]*(-2)+in_buf[767]*(1)+in_buf[768]*(1)+in_buf[769]*(0)+in_buf[770]*(0)+in_buf[771]*(2)+in_buf[772]*(0)+in_buf[773]*(2)+in_buf[774]*(4)+in_buf[775]*(2)+in_buf[776]*(1)+in_buf[777]*(-2)+in_buf[778]*(2)+in_buf[779]*(4)+in_buf[780]*(0)+in_buf[781]*(2)+in_buf[782]*(4)+in_buf[783]*(3);
assign in_buf_weight07=in_buf[0]*(2)+in_buf[1]*(3)+in_buf[2]*(0)+in_buf[3]*(4)+in_buf[4]*(3)+in_buf[5]*(3)+in_buf[6]*(-3)+in_buf[7]*(4)+in_buf[8]*(-3)+in_buf[9]*(-2)+in_buf[10]*(-1)+in_buf[11]*(1)+in_buf[12]*(-7)+in_buf[13]*(-15)+in_buf[14]*(-24)+in_buf[15]*(-16)+in_buf[16]*(3)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(-3)+in_buf[20]*(3)+in_buf[21]*(2)+in_buf[22]*(3)+in_buf[23]*(2)+in_buf[24]*(0)+in_buf[25]*(2)+in_buf[26]*(1)+in_buf[27]*(3)+in_buf[28]*(4)+in_buf[29]*(0)+in_buf[30]*(-3)+in_buf[31]*(1)+in_buf[32]*(0)+in_buf[33]*(-4)+in_buf[34]*(-11)+in_buf[35]*(-11)+in_buf[36]*(-4)+in_buf[37]*(-3)+in_buf[38]*(-10)+in_buf[39]*(-22)+in_buf[40]*(-29)+in_buf[41]*(0)+in_buf[42]*(10)+in_buf[43]*(-43)+in_buf[44]*(-17)+in_buf[45]*(-29)+in_buf[46]*(-28)+in_buf[47]*(-29)+in_buf[48]*(-20)+in_buf[49]*(-14)+in_buf[50]*(-14)+in_buf[51]*(-7)+in_buf[52]*(-2)+in_buf[53]*(0)+in_buf[54]*(2)+in_buf[55]*(-3)+in_buf[56]*(0)+in_buf[57]*(0)+in_buf[58]*(-12)+in_buf[59]*(-31)+in_buf[60]*(-32)+in_buf[61]*(-6)+in_buf[62]*(-6)+in_buf[63]*(-5)+in_buf[64]*(4)+in_buf[65]*(5)+in_buf[66]*(-12)+in_buf[67]*(-18)+in_buf[68]*(-15)+in_buf[69]*(-22)+in_buf[70]*(-2)+in_buf[71]*(-15)+in_buf[72]*(-16)+in_buf[73]*(-15)+in_buf[74]*(-27)+in_buf[75]*(-23)+in_buf[76]*(-22)+in_buf[77]*(-13)+in_buf[78]*(-20)+in_buf[79]*(-22)+in_buf[80]*(0)+in_buf[81]*(-2)+in_buf[82]*(2)+in_buf[83]*(0)+in_buf[84]*(0)+in_buf[85]*(-2)+in_buf[86]*(-16)+in_buf[87]*(-29)+in_buf[88]*(-28)+in_buf[89]*(11)+in_buf[90]*(-8)+in_buf[91]*(14)+in_buf[92]*(3)+in_buf[93]*(-1)+in_buf[94]*(14)+in_buf[95]*(21)+in_buf[96]*(3)+in_buf[97]*(3)+in_buf[98]*(8)+in_buf[99]*(4)+in_buf[100]*(5)+in_buf[101]*(-3)+in_buf[102]*(-16)+in_buf[103]*(-9)+in_buf[104]*(4)+in_buf[105]*(-1)+in_buf[106]*(-7)+in_buf[107]*(-5)+in_buf[108]*(10)+in_buf[109]*(28)+in_buf[110]*(15)+in_buf[111]*(1)+in_buf[112]*(3)+in_buf[113]*(-1)+in_buf[114]*(-28)+in_buf[115]*(1)+in_buf[116]*(0)+in_buf[117]*(-26)+in_buf[118]*(-1)+in_buf[119]*(20)+in_buf[120]*(-18)+in_buf[121]*(2)+in_buf[122]*(6)+in_buf[123]*(12)+in_buf[124]*(3)+in_buf[125]*(-12)+in_buf[126]*(-1)+in_buf[127]*(10)+in_buf[128]*(13)+in_buf[129]*(20)+in_buf[130]*(12)+in_buf[131]*(1)+in_buf[132]*(12)+in_buf[133]*(18)+in_buf[134]*(-1)+in_buf[135]*(8)+in_buf[136]*(33)+in_buf[137]*(30)+in_buf[138]*(-9)+in_buf[139]*(16)+in_buf[140]*(4)+in_buf[141]*(0)+in_buf[142]*(-34)+in_buf[143]*(-6)+in_buf[144]*(-20)+in_buf[145]*(-35)+in_buf[146]*(-14)+in_buf[147]*(-12)+in_buf[148]*(-6)+in_buf[149]*(17)+in_buf[150]*(19)+in_buf[151]*(23)+in_buf[152]*(11)+in_buf[153]*(4)+in_buf[154]*(11)+in_buf[155]*(3)+in_buf[156]*(11)+in_buf[157]*(15)+in_buf[158]*(3)+in_buf[159]*(4)+in_buf[160]*(5)+in_buf[161]*(14)+in_buf[162]*(-13)+in_buf[163]*(-19)+in_buf[164]*(-10)+in_buf[165]*(-8)+in_buf[166]*(10)+in_buf[167]*(13)+in_buf[168]*(2)+in_buf[169]*(-5)+in_buf[170]*(32)+in_buf[171]*(6)+in_buf[172]*(5)+in_buf[173]*(0)+in_buf[174]*(-9)+in_buf[175]*(0)+in_buf[176]*(1)+in_buf[177]*(13)+in_buf[178]*(7)+in_buf[179]*(10)+in_buf[180]*(1)+in_buf[181]*(3)+in_buf[182]*(4)+in_buf[183]*(3)+in_buf[184]*(1)+in_buf[185]*(-2)+in_buf[186]*(-7)+in_buf[187]*(1)+in_buf[188]*(4)+in_buf[189]*(-9)+in_buf[190]*(-10)+in_buf[191]*(11)+in_buf[192]*(6)+in_buf[193]*(-16)+in_buf[194]*(-16)+in_buf[195]*(-12)+in_buf[196]*(-2)+in_buf[197]*(-22)+in_buf[198]*(22)+in_buf[199]*(-6)+in_buf[200]*(-8)+in_buf[201]*(19)+in_buf[202]*(14)+in_buf[203]*(-9)+in_buf[204]*(12)+in_buf[205]*(2)+in_buf[206]*(-4)+in_buf[207]*(1)+in_buf[208]*(-1)+in_buf[209]*(0)+in_buf[210]*(1)+in_buf[211]*(4)+in_buf[212]*(-2)+in_buf[213]*(-1)+in_buf[214]*(-13)+in_buf[215]*(-13)+in_buf[216]*(-8)+in_buf[217]*(-10)+in_buf[218]*(5)+in_buf[219]*(4)+in_buf[220]*(28)+in_buf[221]*(30)+in_buf[222]*(7)+in_buf[223]*(0)+in_buf[224]*(-10)+in_buf[225]*(-13)+in_buf[226]*(17)+in_buf[227]*(0)+in_buf[228]*(-7)+in_buf[229]*(8)+in_buf[230]*(11)+in_buf[231]*(-12)+in_buf[232]*(-7)+in_buf[233]*(-7)+in_buf[234]*(-20)+in_buf[235]*(2)+in_buf[236]*(-6)+in_buf[237]*(-8)+in_buf[238]*(4)+in_buf[239]*(-1)+in_buf[240]*(4)+in_buf[241]*(-3)+in_buf[242]*(-5)+in_buf[243]*(-6)+in_buf[244]*(-6)+in_buf[245]*(11)+in_buf[246]*(-11)+in_buf[247]*(-11)+in_buf[248]*(44)+in_buf[249]*(74)+in_buf[250]*(11)+in_buf[251]*(-1)+in_buf[252]*(-8)+in_buf[253]*(1)+in_buf[254]*(10)+in_buf[255]*(0)+in_buf[256]*(-22)+in_buf[257]*(-14)+in_buf[258]*(8)+in_buf[259]*(-10)+in_buf[260]*(-10)+in_buf[261]*(-6)+in_buf[262]*(-12)+in_buf[263]*(9)+in_buf[264]*(1)+in_buf[265]*(-12)+in_buf[266]*(-19)+in_buf[267]*(-2)+in_buf[268]*(10)+in_buf[269]*(18)+in_buf[270]*(12)+in_buf[271]*(-4)+in_buf[272]*(-4)+in_buf[273]*(-2)+in_buf[274]*(-25)+in_buf[275]*(-13)+in_buf[276]*(24)+in_buf[277]*(19)+in_buf[278]*(21)+in_buf[279]*(-8)+in_buf[280]*(-3)+in_buf[281]*(-4)+in_buf[282]*(-2)+in_buf[283]*(22)+in_buf[284]*(-14)+in_buf[285]*(-1)+in_buf[286]*(1)+in_buf[287]*(0)+in_buf[288]*(0)+in_buf[289]*(0)+in_buf[290]*(0)+in_buf[291]*(4)+in_buf[292]*(-5)+in_buf[293]*(-27)+in_buf[294]*(-23)+in_buf[295]*(-10)+in_buf[296]*(0)+in_buf[297]*(9)+in_buf[298]*(20)+in_buf[299]*(1)+in_buf[300]*(-9)+in_buf[301]*(-14)+in_buf[302]*(-17)+in_buf[303]*(-11)+in_buf[304]*(6)+in_buf[305]*(25)+in_buf[306]*(21)+in_buf[307]*(-9)+in_buf[308]*(-4)+in_buf[309]*(-34)+in_buf[310]*(-32)+in_buf[311]*(-10)+in_buf[312]*(-33)+in_buf[313]*(-5)+in_buf[314]*(16)+in_buf[315]*(-6)+in_buf[316]*(1)+in_buf[317]*(8)+in_buf[318]*(14)+in_buf[319]*(-4)+in_buf[320]*(-14)+in_buf[321]*(-24)+in_buf[322]*(-18)+in_buf[323]*(-5)+in_buf[324]*(7)+in_buf[325]*(13)+in_buf[326]*(7)+in_buf[327]*(5)+in_buf[328]*(-18)+in_buf[329]*(-16)+in_buf[330]*(-19)+in_buf[331]*(-23)+in_buf[332]*(-21)+in_buf[333]*(0)+in_buf[334]*(1)+in_buf[335]*(-2)+in_buf[336]*(-14)+in_buf[337]*(-2)+in_buf[338]*(-8)+in_buf[339]*(-25)+in_buf[340]*(-15)+in_buf[341]*(3)+in_buf[342]*(17)+in_buf[343]*(-2)+in_buf[344]*(-6)+in_buf[345]*(-7)+in_buf[346]*(8)+in_buf[347]*(-7)+in_buf[348]*(-26)+in_buf[349]*(-29)+in_buf[350]*(-17)+in_buf[351]*(-10)+in_buf[352]*(-14)+in_buf[353]*(-1)+in_buf[354]*(3)+in_buf[355]*(6)+in_buf[356]*(-6)+in_buf[357]*(-2)+in_buf[358]*(-13)+in_buf[359]*(-6)+in_buf[360]*(-19)+in_buf[361]*(-2)+in_buf[362]*(12)+in_buf[363]*(-12)+in_buf[364]*(-1)+in_buf[365]*(-4)+in_buf[366]*(-9)+in_buf[367]*(-30)+in_buf[368]*(0)+in_buf[369]*(0)+in_buf[370]*(-5)+in_buf[371]*(14)+in_buf[372]*(9)+in_buf[373]*(15)+in_buf[374]*(22)+in_buf[375]*(-10)+in_buf[376]*(-29)+in_buf[377]*(-26)+in_buf[378]*(-13)+in_buf[379]*(-8)+in_buf[380]*(-12)+in_buf[381]*(-4)+in_buf[382]*(6)+in_buf[383]*(15)+in_buf[384]*(2)+in_buf[385]*(8)+in_buf[386]*(4)+in_buf[387]*(9)+in_buf[388]*(3)+in_buf[389]*(6)+in_buf[390]*(9)+in_buf[391]*(0)+in_buf[392]*(17)+in_buf[393]*(-4)+in_buf[394]*(-23)+in_buf[395]*(-7)+in_buf[396]*(17)+in_buf[397]*(4)+in_buf[398]*(14)+in_buf[399]*(26)+in_buf[400]*(18)+in_buf[401]*(16)+in_buf[402]*(17)+in_buf[403]*(-2)+in_buf[404]*(-22)+in_buf[405]*(-10)+in_buf[406]*(0)+in_buf[407]*(0)+in_buf[408]*(-8)+in_buf[409]*(6)+in_buf[410]*(12)+in_buf[411]*(13)+in_buf[412]*(18)+in_buf[413]*(16)+in_buf[414]*(6)+in_buf[415]*(1)+in_buf[416]*(0)+in_buf[417]*(26)+in_buf[418]*(7)+in_buf[419]*(-8)+in_buf[420]*(9)+in_buf[421]*(1)+in_buf[422]*(-6)+in_buf[423]*(7)+in_buf[424]*(29)+in_buf[425]*(4)+in_buf[426]*(17)+in_buf[427]*(31)+in_buf[428]*(18)+in_buf[429]*(16)+in_buf[430]*(18)+in_buf[431]*(3)+in_buf[432]*(2)+in_buf[433]*(1)+in_buf[434]*(-5)+in_buf[435]*(-2)+in_buf[436]*(-4)+in_buf[437]*(-2)+in_buf[438]*(-2)+in_buf[439]*(18)+in_buf[440]*(7)+in_buf[441]*(6)+in_buf[442]*(2)+in_buf[443]*(9)+in_buf[444]*(-5)+in_buf[445]*(25)+in_buf[446]*(36)+in_buf[447]*(4)+in_buf[448]*(-3)+in_buf[449]*(-12)+in_buf[450]*(0)+in_buf[451]*(24)+in_buf[452]*(11)+in_buf[453]*(26)+in_buf[454]*(30)+in_buf[455]*(28)+in_buf[456]*(26)+in_buf[457]*(0)+in_buf[458]*(7)+in_buf[459]*(18)+in_buf[460]*(24)+in_buf[461]*(12)+in_buf[462]*(-3)+in_buf[463]*(7)+in_buf[464]*(-5)+in_buf[465]*(1)+in_buf[466]*(20)+in_buf[467]*(29)+in_buf[468]*(31)+in_buf[469]*(0)+in_buf[470]*(18)+in_buf[471]*(19)+in_buf[472]*(-6)+in_buf[473]*(38)+in_buf[474]*(28)+in_buf[475]*(-10)+in_buf[476]*(0)+in_buf[477]*(-6)+in_buf[478]*(19)+in_buf[479]*(22)+in_buf[480]*(20)+in_buf[481]*(28)+in_buf[482]*(45)+in_buf[483]*(43)+in_buf[484]*(38)+in_buf[485]*(23)+in_buf[486]*(31)+in_buf[487]*(18)+in_buf[488]*(25)+in_buf[489]*(15)+in_buf[490]*(5)+in_buf[491]*(5)+in_buf[492]*(8)+in_buf[493]*(9)+in_buf[494]*(28)+in_buf[495]*(13)+in_buf[496]*(15)+in_buf[497]*(7)+in_buf[498]*(-8)+in_buf[499]*(-5)+in_buf[500]*(-11)+in_buf[501]*(16)+in_buf[502]*(20)+in_buf[503]*(5)+in_buf[504]*(0)+in_buf[505]*(-11)+in_buf[506]*(0)+in_buf[507]*(14)+in_buf[508]*(30)+in_buf[509]*(24)+in_buf[510]*(45)+in_buf[511]*(45)+in_buf[512]*(24)+in_buf[513]*(26)+in_buf[514]*(31)+in_buf[515]*(35)+in_buf[516]*(38)+in_buf[517]*(33)+in_buf[518]*(2)+in_buf[519]*(-2)+in_buf[520]*(16)+in_buf[521]*(19)+in_buf[522]*(13)+in_buf[523]*(24)+in_buf[524]*(17)+in_buf[525]*(7)+in_buf[526]*(-11)+in_buf[527]*(-6)+in_buf[528]*(-2)+in_buf[529]*(-17)+in_buf[530]*(-12)+in_buf[531]*(-5)+in_buf[532]*(-3)+in_buf[533]*(-7)+in_buf[534]*(6)+in_buf[535]*(22)+in_buf[536]*(25)+in_buf[537]*(15)+in_buf[538]*(19)+in_buf[539]*(15)+in_buf[540]*(17)+in_buf[541]*(7)+in_buf[542]*(19)+in_buf[543]*(31)+in_buf[544]*(21)+in_buf[545]*(4)+in_buf[546]*(8)+in_buf[547]*(5)+in_buf[548]*(10)+in_buf[549]*(16)+in_buf[550]*(33)+in_buf[551]*(22)+in_buf[552]*(13)+in_buf[553]*(10)+in_buf[554]*(-5)+in_buf[555]*(-10)+in_buf[556]*(7)+in_buf[557]*(-12)+in_buf[558]*(43)+in_buf[559]*(1)+in_buf[560]*(-1)+in_buf[561]*(18)+in_buf[562]*(-9)+in_buf[563]*(17)+in_buf[564]*(17)+in_buf[565]*(-1)+in_buf[566]*(-16)+in_buf[567]*(-17)+in_buf[568]*(-8)+in_buf[569]*(-5)+in_buf[570]*(0)+in_buf[571]*(-5)+in_buf[572]*(-16)+in_buf[573]*(-7)+in_buf[574]*(-4)+in_buf[575]*(-2)+in_buf[576]*(7)+in_buf[577]*(18)+in_buf[578]*(14)+in_buf[579]*(16)+in_buf[580]*(13)+in_buf[581]*(8)+in_buf[582]*(0)+in_buf[583]*(-2)+in_buf[584]*(23)+in_buf[585]*(14)+in_buf[586]*(19)+in_buf[587]*(7)+in_buf[588]*(-4)+in_buf[589]*(6)+in_buf[590]*(-28)+in_buf[591]*(-19)+in_buf[592]*(2)+in_buf[593]*(1)+in_buf[594]*(-20)+in_buf[595]*(-21)+in_buf[596]*(-17)+in_buf[597]*(-17)+in_buf[598]*(-24)+in_buf[599]*(-13)+in_buf[600]*(-10)+in_buf[601]*(-10)+in_buf[602]*(4)+in_buf[603]*(15)+in_buf[604]*(23)+in_buf[605]*(15)+in_buf[606]*(12)+in_buf[607]*(6)+in_buf[608]*(17)+in_buf[609]*(13)+in_buf[610]*(17)+in_buf[611]*(26)+in_buf[612]*(30)+in_buf[613]*(-8)+in_buf[614]*(-19)+in_buf[615]*(1)+in_buf[616]*(-3)+in_buf[617]*(9)+in_buf[618]*(-10)+in_buf[619]*(-26)+in_buf[620]*(-6)+in_buf[621]*(-22)+in_buf[622]*(-30)+in_buf[623]*(-34)+in_buf[624]*(-27)+in_buf[625]*(-33)+in_buf[626]*(-26)+in_buf[627]*(-7)+in_buf[628]*(-2)+in_buf[629]*(-3)+in_buf[630]*(19)+in_buf[631]*(22)+in_buf[632]*(28)+in_buf[633]*(19)+in_buf[634]*(2)+in_buf[635]*(6)+in_buf[636]*(6)+in_buf[637]*(21)+in_buf[638]*(31)+in_buf[639]*(45)+in_buf[640]*(41)+in_buf[641]*(-3)+in_buf[642]*(-5)+in_buf[643]*(3)+in_buf[644]*(3)+in_buf[645]*(-2)+in_buf[646]*(-4)+in_buf[647]*(10)+in_buf[648]*(-10)+in_buf[649]*(-11)+in_buf[650]*(-21)+in_buf[651]*(-15)+in_buf[652]*(-4)+in_buf[653]*(-21)+in_buf[654]*(-16)+in_buf[655]*(0)+in_buf[656]*(-11)+in_buf[657]*(5)+in_buf[658]*(24)+in_buf[659]*(32)+in_buf[660]*(25)+in_buf[661]*(10)+in_buf[662]*(9)+in_buf[663]*(1)+in_buf[664]*(20)+in_buf[665]*(44)+in_buf[666]*(20)+in_buf[667]*(36)+in_buf[668]*(38)+in_buf[669]*(5)+in_buf[670]*(1)+in_buf[671]*(4)+in_buf[672]*(0)+in_buf[673]*(2)+in_buf[674]*(-14)+in_buf[675]*(4)+in_buf[676]*(-1)+in_buf[677]*(-15)+in_buf[678]*(-11)+in_buf[679]*(3)+in_buf[680]*(1)+in_buf[681]*(4)+in_buf[682]*(1)+in_buf[683]*(7)+in_buf[684]*(4)+in_buf[685]*(5)+in_buf[686]*(17)+in_buf[687]*(22)+in_buf[688]*(26)+in_buf[689]*(8)+in_buf[690]*(-4)+in_buf[691]*(-7)+in_buf[692]*(31)+in_buf[693]*(31)+in_buf[694]*(42)+in_buf[695]*(56)+in_buf[696]*(-7)+in_buf[697]*(17)+in_buf[698]*(5)+in_buf[699]*(-3)+in_buf[700]*(0)+in_buf[701]*(-3)+in_buf[702]*(31)+in_buf[703]*(6)+in_buf[704]*(-6)+in_buf[705]*(-5)+in_buf[706]*(15)+in_buf[707]*(4)+in_buf[708]*(-1)+in_buf[709]*(-11)+in_buf[710]*(8)+in_buf[711]*(18)+in_buf[712]*(-17)+in_buf[713]*(-5)+in_buf[714]*(4)+in_buf[715]*(16)+in_buf[716]*(3)+in_buf[717]*(-12)+in_buf[718]*(0)+in_buf[719]*(5)+in_buf[720]*(19)+in_buf[721]*(26)+in_buf[722]*(38)+in_buf[723]*(22)+in_buf[724]*(-11)+in_buf[725]*(22)+in_buf[726]*(3)+in_buf[727]*(1)+in_buf[728]*(2)+in_buf[729]*(3)+in_buf[730]*(0)+in_buf[731]*(0)+in_buf[732]*(19)+in_buf[733]*(18)+in_buf[734]*(28)+in_buf[735]*(0)+in_buf[736]*(24)+in_buf[737]*(0)+in_buf[738]*(10)+in_buf[739]*(6)+in_buf[740]*(38)+in_buf[741]*(20)+in_buf[742]*(5)+in_buf[743]*(14)+in_buf[744]*(-6)+in_buf[745]*(-12)+in_buf[746]*(-15)+in_buf[747]*(-17)+in_buf[748]*(-5)+in_buf[749]*(2)+in_buf[750]*(8)+in_buf[751]*(27)+in_buf[752]*(23)+in_buf[753]*(-4)+in_buf[754]*(0)+in_buf[755]*(3)+in_buf[756]*(-3)+in_buf[757]*(0)+in_buf[758]*(-1)+in_buf[759]*(0)+in_buf[760]*(-4)+in_buf[761]*(0)+in_buf[762]*(1)+in_buf[763]*(8)+in_buf[764]*(3)+in_buf[765]*(-7)+in_buf[766]*(6)+in_buf[767]*(2)+in_buf[768]*(-1)+in_buf[769]*(-37)+in_buf[770]*(-23)+in_buf[771]*(3)+in_buf[772]*(-26)+in_buf[773]*(-42)+in_buf[774]*(-25)+in_buf[775]*(21)+in_buf[776]*(13)+in_buf[777]*(-14)+in_buf[778]*(-6)+in_buf[779]*(-22)+in_buf[780]*(-2)+in_buf[781]*(0)+in_buf[782]*(2)+in_buf[783]*(-1);
assign in_buf_weight08=in_buf[0]*(4)+in_buf[1]*(-3)+in_buf[2]*(2)+in_buf[3]*(0)+in_buf[4]*(-1)+in_buf[5]*(0)+in_buf[6]*(-2)+in_buf[7]*(-1)+in_buf[8]*(-4)+in_buf[9]*(0)+in_buf[10]*(3)+in_buf[11]*(3)+in_buf[12]*(5)+in_buf[13]*(3)+in_buf[14]*(4)+in_buf[15]*(3)+in_buf[16]*(-3)+in_buf[17]*(-2)+in_buf[18]*(3)+in_buf[19]*(-2)+in_buf[20]*(-2)+in_buf[21]*(2)+in_buf[22]*(2)+in_buf[23]*(-2)+in_buf[24]*(-3)+in_buf[25]*(-1)+in_buf[26]*(3)+in_buf[27]*(-1)+in_buf[28]*(0)+in_buf[29]*(2)+in_buf[30]*(4)+in_buf[31]*(-3)+in_buf[32]*(5)+in_buf[33]*(2)+in_buf[34]*(0)+in_buf[35]*(9)+in_buf[36]*(2)+in_buf[37]*(9)+in_buf[38]*(3)+in_buf[39]*(13)+in_buf[40]*(21)+in_buf[41]*(14)+in_buf[42]*(19)+in_buf[43]*(34)+in_buf[44]*(12)+in_buf[45]*(14)+in_buf[46]*(10)+in_buf[47]*(16)+in_buf[48]*(6)+in_buf[49]*(10)+in_buf[50]*(8)+in_buf[51]*(8)+in_buf[52]*(2)+in_buf[53]*(-1)+in_buf[54]*(-2)+in_buf[55]*(-1)+in_buf[56]*(-1)+in_buf[57]*(4)+in_buf[58]*(2)+in_buf[59]*(23)+in_buf[60]*(35)+in_buf[61]*(1)+in_buf[62]*(2)+in_buf[63]*(19)+in_buf[64]*(6)+in_buf[65]*(5)+in_buf[66]*(28)+in_buf[67]*(27)+in_buf[68]*(27)+in_buf[69]*(28)+in_buf[70]*(6)+in_buf[71]*(0)+in_buf[72]*(20)+in_buf[73]*(36)+in_buf[74]*(45)+in_buf[75]*(30)+in_buf[76]*(17)+in_buf[77]*(12)+in_buf[78]*(24)+in_buf[79]*(14)+in_buf[80]*(-2)+in_buf[81]*(-2)+in_buf[82]*(0)+in_buf[83]*(2)+in_buf[84]*(-3)+in_buf[85]*(-3)+in_buf[86]*(22)+in_buf[87]*(33)+in_buf[88]*(30)+in_buf[89]*(-11)+in_buf[90]*(-18)+in_buf[91]*(2)+in_buf[92]*(10)+in_buf[93]*(-18)+in_buf[94]*(-6)+in_buf[95]*(-16)+in_buf[96]*(3)+in_buf[97]*(16)+in_buf[98]*(29)+in_buf[99]*(24)+in_buf[100]*(17)+in_buf[101]*(20)+in_buf[102]*(20)+in_buf[103]*(0)+in_buf[104]*(-24)+in_buf[105]*(-18)+in_buf[106]*(4)+in_buf[107]*(22)+in_buf[108]*(0)+in_buf[109]*(-14)+in_buf[110]*(-24)+in_buf[111]*(-1)+in_buf[112]*(4)+in_buf[113]*(1)+in_buf[114]*(16)+in_buf[115]*(9)+in_buf[116]*(-8)+in_buf[117]*(-17)+in_buf[118]*(-13)+in_buf[119]*(6)+in_buf[120]*(13)+in_buf[121]*(-2)+in_buf[122]*(-17)+in_buf[123]*(-18)+in_buf[124]*(-10)+in_buf[125]*(-7)+in_buf[126]*(13)+in_buf[127]*(33)+in_buf[128]*(20)+in_buf[129]*(11)+in_buf[130]*(3)+in_buf[131]*(7)+in_buf[132]*(-20)+in_buf[133]*(-18)+in_buf[134]*(0)+in_buf[135]*(-17)+in_buf[136]*(-46)+in_buf[137]*(-9)+in_buf[138]*(30)+in_buf[139]*(8)+in_buf[140]*(3)+in_buf[141]*(-2)+in_buf[142]*(18)+in_buf[143]*(3)+in_buf[144]*(-18)+in_buf[145]*(-25)+in_buf[146]*(-10)+in_buf[147]*(0)+in_buf[148]*(8)+in_buf[149]*(-11)+in_buf[150]*(-14)+in_buf[151]*(-26)+in_buf[152]*(-23)+in_buf[153]*(5)+in_buf[154]*(15)+in_buf[155]*(15)+in_buf[156]*(0)+in_buf[157]*(7)+in_buf[158]*(12)+in_buf[159]*(5)+in_buf[160]*(-3)+in_buf[161]*(7)+in_buf[162]*(-3)+in_buf[163]*(-37)+in_buf[164]*(-27)+in_buf[165]*(-11)+in_buf[166]*(-2)+in_buf[167]*(-16)+in_buf[168]*(-2)+in_buf[169]*(15)+in_buf[170]*(-7)+in_buf[171]*(15)+in_buf[172]*(-25)+in_buf[173]*(-20)+in_buf[174]*(8)+in_buf[175]*(4)+in_buf[176]*(-5)+in_buf[177]*(-32)+in_buf[178]*(-21)+in_buf[179]*(-32)+in_buf[180]*(-15)+in_buf[181]*(-4)+in_buf[182]*(3)+in_buf[183]*(1)+in_buf[184]*(4)+in_buf[185]*(16)+in_buf[186]*(29)+in_buf[187]*(10)+in_buf[188]*(16)+in_buf[189]*(19)+in_buf[190]*(-5)+in_buf[191]*(-22)+in_buf[192]*(-21)+in_buf[193]*(-14)+in_buf[194]*(-7)+in_buf[195]*(-17)+in_buf[196]*(-2)+in_buf[197]*(3)+in_buf[198]*(-13)+in_buf[199]*(17)+in_buf[200]*(-9)+in_buf[201]*(-22)+in_buf[202]*(-19)+in_buf[203]*(-16)+in_buf[204]*(-18)+in_buf[205]*(-37)+in_buf[206]*(-25)+in_buf[207]*(-11)+in_buf[208]*(-6)+in_buf[209]*(-6)+in_buf[210]*(4)+in_buf[211]*(21)+in_buf[212]*(29)+in_buf[213]*(31)+in_buf[214]*(39)+in_buf[215]*(28)+in_buf[216]*(25)+in_buf[217]*(30)+in_buf[218]*(15)+in_buf[219]*(0)+in_buf[220]*(-16)+in_buf[221]*(-10)+in_buf[222]*(-9)+in_buf[223]*(-15)+in_buf[224]*(34)+in_buf[225]*(-5)+in_buf[226]*(-17)+in_buf[227]*(-8)+in_buf[228]*(-19)+in_buf[229]*(-14)+in_buf[230]*(-2)+in_buf[231]*(-4)+in_buf[232]*(-8)+in_buf[233]*(-27)+in_buf[234]*(-13)+in_buf[235]*(-14)+in_buf[236]*(-3)+in_buf[237]*(0)+in_buf[238]*(20)+in_buf[239]*(24)+in_buf[240]*(43)+in_buf[241]*(39)+in_buf[242]*(24)+in_buf[243]*(26)+in_buf[244]*(28)+in_buf[245]*(26)+in_buf[246]*(28)+in_buf[247]*(5)+in_buf[248]*(-4)+in_buf[249]*(-10)+in_buf[250]*(-5)+in_buf[251]*(15)+in_buf[252]*(6)+in_buf[253]*(19)+in_buf[254]*(-20)+in_buf[255]*(-2)+in_buf[256]*(-16)+in_buf[257]*(-21)+in_buf[258]*(-6)+in_buf[259]*(0)+in_buf[260]*(11)+in_buf[261]*(1)+in_buf[262]*(3)+in_buf[263]*(-23)+in_buf[264]*(0)+in_buf[265]*(9)+in_buf[266]*(4)+in_buf[267]*(18)+in_buf[268]*(27)+in_buf[269]*(12)+in_buf[270]*(2)+in_buf[271]*(17)+in_buf[272]*(24)+in_buf[273]*(15)+in_buf[274]*(18)+in_buf[275]*(14)+in_buf[276]*(10)+in_buf[277]*(35)+in_buf[278]*(11)+in_buf[279]*(13)+in_buf[280]*(10)+in_buf[281]*(15)+in_buf[282]*(1)+in_buf[283]*(-3)+in_buf[284]*(-28)+in_buf[285]*(-12)+in_buf[286]*(-3)+in_buf[287]*(9)+in_buf[288]*(11)+in_buf[289]*(0)+in_buf[290]*(1)+in_buf[291]*(-3)+in_buf[292]*(-1)+in_buf[293]*(1)+in_buf[294]*(6)+in_buf[295]*(18)+in_buf[296]*(15)+in_buf[297]*(-5)+in_buf[298]*(7)+in_buf[299]*(4)+in_buf[300]*(22)+in_buf[301]*(16)+in_buf[302]*(29)+in_buf[303]*(39)+in_buf[304]*(29)+in_buf[305]*(16)+in_buf[306]*(30)+in_buf[307]*(14)+in_buf[308]*(8)+in_buf[309]*(13)+in_buf[310]*(7)+in_buf[311]*(-11)+in_buf[312]*(-13)+in_buf[313]*(-7)+in_buf[314]*(-1)+in_buf[315]*(23)+in_buf[316]*(6)+in_buf[317]*(-2)+in_buf[318]*(9)+in_buf[319]*(25)+in_buf[320]*(-7)+in_buf[321]*(-2)+in_buf[322]*(3)+in_buf[323]*(-3)+in_buf[324]*(-17)+in_buf[325]*(-9)+in_buf[326]*(4)+in_buf[327]*(-6)+in_buf[328]*(23)+in_buf[329]*(37)+in_buf[330]*(38)+in_buf[331]*(44)+in_buf[332]*(52)+in_buf[333]*(37)+in_buf[334]*(66)+in_buf[335]*(38)+in_buf[336]*(14)+in_buf[337]*(5)+in_buf[338]*(16)+in_buf[339]*(-2)+in_buf[340]*(12)+in_buf[341]*(17)+in_buf[342]*(25)+in_buf[343]*(13)+in_buf[344]*(3)+in_buf[345]*(9)+in_buf[346]*(8)+in_buf[347]*(11)+in_buf[348]*(-34)+in_buf[349]*(-43)+in_buf[350]*(-6)+in_buf[351]*(-14)+in_buf[352]*(-26)+in_buf[353]*(-16)+in_buf[354]*(-16)+in_buf[355]*(-12)+in_buf[356]*(9)+in_buf[357]*(20)+in_buf[358]*(25)+in_buf[359]*(37)+in_buf[360]*(26)+in_buf[361]*(15)+in_buf[362]*(30)+in_buf[363]*(38)+in_buf[364]*(22)+in_buf[365]*(10)+in_buf[366]*(17)+in_buf[367]*(-6)+in_buf[368]*(2)+in_buf[369]*(5)+in_buf[370]*(16)+in_buf[371]*(-8)+in_buf[372]*(-5)+in_buf[373]*(-7)+in_buf[374]*(2)+in_buf[375]*(5)+in_buf[376]*(-14)+in_buf[377]*(-23)+in_buf[378]*(-1)+in_buf[379]*(-10)+in_buf[380]*(-22)+in_buf[381]*(-23)+in_buf[382]*(-30)+in_buf[383]*(-20)+in_buf[384]*(-5)+in_buf[385]*(3)+in_buf[386]*(7)+in_buf[387]*(13)+in_buf[388]*(-12)+in_buf[389]*(1)+in_buf[390]*(8)+in_buf[391]*(10)+in_buf[392]*(11)+in_buf[393]*(6)+in_buf[394]*(25)+in_buf[395]*(-3)+in_buf[396]*(-13)+in_buf[397]*(4)+in_buf[398]*(5)+in_buf[399]*(-21)+in_buf[400]*(-17)+in_buf[401]*(-8)+in_buf[402]*(1)+in_buf[403]*(12)+in_buf[404]*(-4)+in_buf[405]*(1)+in_buf[406]*(6)+in_buf[407]*(2)+in_buf[408]*(-19)+in_buf[409]*(-23)+in_buf[410]*(-26)+in_buf[411]*(-24)+in_buf[412]*(4)+in_buf[413]*(17)+in_buf[414]*(17)+in_buf[415]*(-5)+in_buf[416]*(-15)+in_buf[417]*(-5)+in_buf[418]*(8)+in_buf[419]*(5)+in_buf[420]*(15)+in_buf[421]*(7)+in_buf[422]*(-3)+in_buf[423]*(-45)+in_buf[424]*(-26)+in_buf[425]*(3)+in_buf[426]*(-4)+in_buf[427]*(-1)+in_buf[428]*(-3)+in_buf[429]*(-8)+in_buf[430]*(-3)+in_buf[431]*(10)+in_buf[432]*(10)+in_buf[433]*(-2)+in_buf[434]*(1)+in_buf[435]*(-9)+in_buf[436]*(-16)+in_buf[437]*(-30)+in_buf[438]*(-17)+in_buf[439]*(-22)+in_buf[440]*(10)+in_buf[441]*(8)+in_buf[442]*(-4)+in_buf[443]*(-26)+in_buf[444]*(-2)+in_buf[445]*(-14)+in_buf[446]*(-19)+in_buf[447]*(-19)+in_buf[448]*(0)+in_buf[449]*(8)+in_buf[450]*(5)+in_buf[451]*(-50)+in_buf[452]*(-34)+in_buf[453]*(-3)+in_buf[454]*(-4)+in_buf[455]*(-8)+in_buf[456]*(2)+in_buf[457]*(9)+in_buf[458]*(13)+in_buf[459]*(8)+in_buf[460]*(-4)+in_buf[461]*(-5)+in_buf[462]*(-18)+in_buf[463]*(-20)+in_buf[464]*(-6)+in_buf[465]*(-25)+in_buf[466]*(-17)+in_buf[467]*(-36)+in_buf[468]*(-28)+in_buf[469]*(-41)+in_buf[470]*(-25)+in_buf[471]*(-23)+in_buf[472]*(14)+in_buf[473]*(-6)+in_buf[474]*(-20)+in_buf[475]*(-16)+in_buf[476]*(0)+in_buf[477]*(12)+in_buf[478]*(-29)+in_buf[479]*(-41)+in_buf[480]*(-31)+in_buf[481]*(-8)+in_buf[482]*(-8)+in_buf[483]*(1)+in_buf[484]*(-8)+in_buf[485]*(-3)+in_buf[486]*(5)+in_buf[487]*(-3)+in_buf[488]*(-10)+in_buf[489]*(-7)+in_buf[490]*(-19)+in_buf[491]*(-20)+in_buf[492]*(-10)+in_buf[493]*(-6)+in_buf[494]*(-10)+in_buf[495]*(-3)+in_buf[496]*(-21)+in_buf[497]*(-44)+in_buf[498]*(-24)+in_buf[499]*(-13)+in_buf[500]*(5)+in_buf[501]*(14)+in_buf[502]*(-22)+in_buf[503]*(-1)+in_buf[504]*(16)+in_buf[505]*(8)+in_buf[506]*(-14)+in_buf[507]*(-45)+in_buf[508]*(-21)+in_buf[509]*(-16)+in_buf[510]*(-7)+in_buf[511]*(17)+in_buf[512]*(1)+in_buf[513]*(6)+in_buf[514]*(6)+in_buf[515]*(-2)+in_buf[516]*(-10)+in_buf[517]*(-12)+in_buf[518]*(-26)+in_buf[519]*(-10)+in_buf[520]*(-19)+in_buf[521]*(7)+in_buf[522]*(3)+in_buf[523]*(-7)+in_buf[524]*(-17)+in_buf[525]*(-7)+in_buf[526]*(2)+in_buf[527]*(-10)+in_buf[528]*(-7)+in_buf[529]*(8)+in_buf[530]*(-27)+in_buf[531]*(-20)+in_buf[532]*(6)+in_buf[533]*(27)+in_buf[534]*(16)+in_buf[535]*(-40)+in_buf[536]*(-8)+in_buf[537]*(-4)+in_buf[538]*(5)+in_buf[539]*(1)+in_buf[540]*(1)+in_buf[541]*(-2)+in_buf[542]*(2)+in_buf[543]*(-8)+in_buf[544]*(10)+in_buf[545]*(-3)+in_buf[546]*(-18)+in_buf[547]*(-6)+in_buf[548]*(-8)+in_buf[549]*(2)+in_buf[550]*(0)+in_buf[551]*(-4)+in_buf[552]*(-1)+in_buf[553]*(1)+in_buf[554]*(16)+in_buf[555]*(-4)+in_buf[556]*(23)+in_buf[557]*(3)+in_buf[558]*(-23)+in_buf[559]*(-15)+in_buf[560]*(1)+in_buf[561]*(27)+in_buf[562]*(20)+in_buf[563]*(-34)+in_buf[564]*(-4)+in_buf[565]*(1)+in_buf[566]*(-6)+in_buf[567]*(-4)+in_buf[568]*(4)+in_buf[569]*(2)+in_buf[570]*(6)+in_buf[571]*(16)+in_buf[572]*(35)+in_buf[573]*(19)+in_buf[574]*(8)+in_buf[575]*(7)+in_buf[576]*(-3)+in_buf[577]*(4)+in_buf[578]*(2)+in_buf[579]*(-1)+in_buf[580]*(1)+in_buf[581]*(18)+in_buf[582]*(19)+in_buf[583]*(2)+in_buf[584]*(24)+in_buf[585]*(18)+in_buf[586]*(-1)+in_buf[587]*(6)+in_buf[588]*(0)+in_buf[589]*(-10)+in_buf[590]*(10)+in_buf[591]*(2)+in_buf[592]*(-8)+in_buf[593]*(-8)+in_buf[594]*(17)+in_buf[595]*(17)+in_buf[596]*(-2)+in_buf[597]*(4)+in_buf[598]*(14)+in_buf[599]*(11)+in_buf[600]*(32)+in_buf[601]*(17)+in_buf[602]*(21)+in_buf[603]*(15)+in_buf[604]*(4)+in_buf[605]*(16)+in_buf[606]*(17)+in_buf[607]*(27)+in_buf[608]*(9)+in_buf[609]*(7)+in_buf[610]*(-5)+in_buf[611]*(0)+in_buf[612]*(12)+in_buf[613]*(18)+in_buf[614]*(23)+in_buf[615]*(6)+in_buf[616]*(4)+in_buf[617]*(0)+in_buf[618]*(6)+in_buf[619]*(-4)+in_buf[620]*(-6)+in_buf[621]*(21)+in_buf[622]*(27)+in_buf[623]*(10)+in_buf[624]*(15)+in_buf[625]*(25)+in_buf[626]*(5)+in_buf[627]*(2)+in_buf[628]*(19)+in_buf[629]*(25)+in_buf[630]*(32)+in_buf[631]*(29)+in_buf[632]*(19)+in_buf[633]*(13)+in_buf[634]*(13)+in_buf[635]*(8)+in_buf[636]*(4)+in_buf[637]*(-21)+in_buf[638]*(-34)+in_buf[639]*(-13)+in_buf[640]*(-10)+in_buf[641]*(17)+in_buf[642]*(15)+in_buf[643]*(3)+in_buf[644]*(1)+in_buf[645]*(1)+in_buf[646]*(21)+in_buf[647]*(-31)+in_buf[648]*(-11)+in_buf[649]*(10)+in_buf[650]*(0)+in_buf[651]*(-7)+in_buf[652]*(-7)+in_buf[653]*(14)+in_buf[654]*(-2)+in_buf[655]*(5)+in_buf[656]*(24)+in_buf[657]*(24)+in_buf[658]*(18)+in_buf[659]*(33)+in_buf[660]*(18)+in_buf[661]*(7)+in_buf[662]*(-19)+in_buf[663]*(-12)+in_buf[664]*(-9)+in_buf[665]*(-29)+in_buf[666]*(-16)+in_buf[667]*(-15)+in_buf[668]*(-16)+in_buf[669]*(-6)+in_buf[670]*(-1)+in_buf[671]*(-3)+in_buf[672]*(2)+in_buf[673]*(-3)+in_buf[674]*(-6)+in_buf[675]*(-15)+in_buf[676]*(18)+in_buf[677]*(17)+in_buf[678]*(-24)+in_buf[679]*(-32)+in_buf[680]*(-9)+in_buf[681]*(0)+in_buf[682]*(9)+in_buf[683]*(0)+in_buf[684]*(14)+in_buf[685]*(15)+in_buf[686]*(4)+in_buf[687]*(26)+in_buf[688]*(8)+in_buf[689]*(8)+in_buf[690]*(-16)+in_buf[691]*(-11)+in_buf[692]*(-14)+in_buf[693]*(-20)+in_buf[694]*(-25)+in_buf[695]*(-24)+in_buf[696]*(-16)+in_buf[697]*(-24)+in_buf[698]*(-4)+in_buf[699]*(0)+in_buf[700]*(4)+in_buf[701]*(3)+in_buf[702]*(-29)+in_buf[703]*(15)+in_buf[704]*(2)+in_buf[705]*(-5)+in_buf[706]*(-13)+in_buf[707]*(-1)+in_buf[708]*(15)+in_buf[709]*(34)+in_buf[710]*(13)+in_buf[711]*(-10)+in_buf[712]*(-1)+in_buf[713]*(1)+in_buf[714]*(5)+in_buf[715]*(0)+in_buf[716]*(6)+in_buf[717]*(-3)+in_buf[718]*(5)+in_buf[719]*(31)+in_buf[720]*(14)+in_buf[721]*(9)+in_buf[722]*(-12)+in_buf[723]*(-18)+in_buf[724]*(-17)+in_buf[725]*(-13)+in_buf[726]*(-3)+in_buf[727]*(-1)+in_buf[728]*(4)+in_buf[729]*(-2)+in_buf[730]*(2)+in_buf[731]*(9)+in_buf[732]*(-18)+in_buf[733]*(-18)+in_buf[734]*(-19)+in_buf[735]*(8)+in_buf[736]*(45)+in_buf[737]*(61)+in_buf[738]*(24)+in_buf[739]*(0)+in_buf[740]*(30)+in_buf[741]*(49)+in_buf[742]*(39)+in_buf[743]*(5)+in_buf[744]*(20)+in_buf[745]*(24)+in_buf[746]*(29)+in_buf[747]*(36)+in_buf[748]*(32)+in_buf[749]*(29)+in_buf[750]*(12)+in_buf[751]*(15)+in_buf[752]*(0)+in_buf[753]*(10)+in_buf[754]*(4)+in_buf[755]*(-3)+in_buf[756]*(2)+in_buf[757]*(3)+in_buf[758]*(4)+in_buf[759]*(-2)+in_buf[760]*(20)+in_buf[761]*(18)+in_buf[762]*(18)+in_buf[763]*(20)+in_buf[764]*(19)+in_buf[765]*(23)+in_buf[766]*(55)+in_buf[767]*(50)+in_buf[768]*(42)+in_buf[769]*(51)+in_buf[770]*(64)+in_buf[771]*(31)+in_buf[772]*(11)+in_buf[773]*(27)+in_buf[774]*(14)+in_buf[775]*(18)+in_buf[776]*(-7)+in_buf[777]*(-5)+in_buf[778]*(-8)+in_buf[779]*(-16)+in_buf[780]*(2)+in_buf[781]*(-1)+in_buf[782]*(1)+in_buf[783]*(2);
assign in_buf_weight09=in_buf[0]*(-3)+in_buf[1]*(0)+in_buf[2]*(0)+in_buf[3]*(-3)+in_buf[4]*(-1)+in_buf[5]*(4)+in_buf[6]*(4)+in_buf[7]*(2)+in_buf[8]*(0)+in_buf[9]*(-3)+in_buf[10]*(1)+in_buf[11]*(-3)+in_buf[12]*(0)+in_buf[13]*(-3)+in_buf[14]*(4)+in_buf[15]*(0)+in_buf[16]*(-2)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(0)+in_buf[20]*(0)+in_buf[21]*(3)+in_buf[22]*(0)+in_buf[23]*(1)+in_buf[24]*(2)+in_buf[25]*(3)+in_buf[26]*(3)+in_buf[27]*(-2)+in_buf[28]*(3)+in_buf[29]*(4)+in_buf[30]*(-3)+in_buf[31]*(-1)+in_buf[32]*(2)+in_buf[33]*(0)+in_buf[34]*(0)+in_buf[35]*(1)+in_buf[36]*(0)+in_buf[37]*(0)+in_buf[38]*(4)+in_buf[39]*(-1)+in_buf[40]*(-2)+in_buf[41]*(1)+in_buf[42]*(-1)+in_buf[43]*(1)+in_buf[44]*(2)+in_buf[45]*(-2)+in_buf[46]*(0)+in_buf[47]*(0)+in_buf[48]*(0)+in_buf[49]*(0)+in_buf[50]*(-1)+in_buf[51]*(-3)+in_buf[52]*(4)+in_buf[53]*(0)+in_buf[54]*(0)+in_buf[55]*(-1)+in_buf[56]*(0)+in_buf[57]*(1)+in_buf[58]*(-2)+in_buf[59]*(1)+in_buf[60]*(1)+in_buf[61]*(3)+in_buf[62]*(4)+in_buf[63]*(-1)+in_buf[64]*(-1)+in_buf[65]*(5)+in_buf[66]*(-1)+in_buf[67]*(-2)+in_buf[68]*(1)+in_buf[69]*(4)+in_buf[70]*(2)+in_buf[71]*(3)+in_buf[72]*(0)+in_buf[73]*(-1)+in_buf[74]*(-2)+in_buf[75]*(-3)+in_buf[76]*(0)+in_buf[77]*(0)+in_buf[78]*(-1)+in_buf[79]*(0)+in_buf[80]*(0)+in_buf[81]*(1)+in_buf[82]*(0)+in_buf[83]*(-1)+in_buf[84]*(0)+in_buf[85]*(0)+in_buf[86]*(4)+in_buf[87]*(-1)+in_buf[88]*(-3)+in_buf[89]*(0)+in_buf[90]*(5)+in_buf[91]*(-2)+in_buf[92]*(-1)+in_buf[93]*(2)+in_buf[94]*(-2)+in_buf[95]*(-1)+in_buf[96]*(0)+in_buf[97]*(6)+in_buf[98]*(4)+in_buf[99]*(1)+in_buf[100]*(0)+in_buf[101]*(-1)+in_buf[102]*(3)+in_buf[103]*(2)+in_buf[104]*(2)+in_buf[105]*(-3)+in_buf[106]*(2)+in_buf[107]*(1)+in_buf[108]*(3)+in_buf[109]*(0)+in_buf[110]*(0)+in_buf[111]*(2)+in_buf[112]*(4)+in_buf[113]*(0)+in_buf[114]*(0)+in_buf[115]*(-5)+in_buf[116]*(0)+in_buf[117]*(2)+in_buf[118]*(-1)+in_buf[119]*(1)+in_buf[120]*(2)+in_buf[121]*(0)+in_buf[122]*(2)+in_buf[123]*(-2)+in_buf[124]*(0)+in_buf[125]*(1)+in_buf[126]*(0)+in_buf[127]*(-2)+in_buf[128]*(-1)+in_buf[129]*(-4)+in_buf[130]*(-4)+in_buf[131]*(0)+in_buf[132]*(0)+in_buf[133]*(2)+in_buf[134]*(-1)+in_buf[135]*(0)+in_buf[136]*(6)+in_buf[137]*(-1)+in_buf[138]*(1)+in_buf[139]*(2)+in_buf[140]*(0)+in_buf[141]*(0)+in_buf[142]*(3)+in_buf[143]*(-3)+in_buf[144]*(-3)+in_buf[145]*(4)+in_buf[146]*(6)+in_buf[147]*(0)+in_buf[148]*(3)+in_buf[149]*(7)+in_buf[150]*(1)+in_buf[151]*(0)+in_buf[152]*(-1)+in_buf[153]*(2)+in_buf[154]*(1)+in_buf[155]*(3)+in_buf[156]*(-2)+in_buf[157]*(0)+in_buf[158]*(0)+in_buf[159]*(0)+in_buf[160]*(-5)+in_buf[161]*(-2)+in_buf[162]*(-3)+in_buf[163]*(0)+in_buf[164]*(5)+in_buf[165]*(5)+in_buf[166]*(4)+in_buf[167]*(3)+in_buf[168]*(-1)+in_buf[169]*(-2)+in_buf[170]*(1)+in_buf[171]*(-2)+in_buf[172]*(-2)+in_buf[173]*(3)+in_buf[174]*(1)+in_buf[175]*(6)+in_buf[176]*(6)+in_buf[177]*(1)+in_buf[178]*(0)+in_buf[179]*(0)+in_buf[180]*(4)+in_buf[181]*(-1)+in_buf[182]*(1)+in_buf[183]*(1)+in_buf[184]*(2)+in_buf[185]*(-2)+in_buf[186]*(0)+in_buf[187]*(-4)+in_buf[188]*(-3)+in_buf[189]*(1)+in_buf[190]*(-1)+in_buf[191]*(4)+in_buf[192]*(0)+in_buf[193]*(-1)+in_buf[194]*(4)+in_buf[195]*(0)+in_buf[196]*(3)+in_buf[197]*(2)+in_buf[198]*(3)+in_buf[199]*(2)+in_buf[200]*(-6)+in_buf[201]*(0)+in_buf[202]*(0)+in_buf[203]*(2)+in_buf[204]*(0)+in_buf[205]*(-4)+in_buf[206]*(3)+in_buf[207]*(-3)+in_buf[208]*(-1)+in_buf[209]*(-3)+in_buf[210]*(-2)+in_buf[211]*(1)+in_buf[212]*(-4)+in_buf[213]*(0)+in_buf[214]*(2)+in_buf[215]*(-1)+in_buf[216]*(-2)+in_buf[217]*(-1)+in_buf[218]*(-2)+in_buf[219]*(0)+in_buf[220]*(0)+in_buf[221]*(0)+in_buf[222]*(-2)+in_buf[223]*(2)+in_buf[224]*(4)+in_buf[225]*(4)+in_buf[226]*(0)+in_buf[227]*(0)+in_buf[228]*(-3)+in_buf[229]*(1)+in_buf[230]*(-2)+in_buf[231]*(0)+in_buf[232]*(-2)+in_buf[233]*(-3)+in_buf[234]*(-1)+in_buf[235]*(-2)+in_buf[236]*(-6)+in_buf[237]*(-4)+in_buf[238]*(-6)+in_buf[239]*(-3)+in_buf[240]*(0)+in_buf[241]*(3)+in_buf[242]*(2)+in_buf[243]*(-4)+in_buf[244]*(-1)+in_buf[245]*(0)+in_buf[246]*(-3)+in_buf[247]*(-3)+in_buf[248]*(6)+in_buf[249]*(3)+in_buf[250]*(2)+in_buf[251]*(0)+in_buf[252]*(4)+in_buf[253]*(0)+in_buf[254]*(-1)+in_buf[255]*(0)+in_buf[256]*(-3)+in_buf[257]*(-3)+in_buf[258]*(-5)+in_buf[259]*(-3)+in_buf[260]*(-2)+in_buf[261]*(-1)+in_buf[262]*(2)+in_buf[263]*(-5)+in_buf[264]*(-3)+in_buf[265]*(-3)+in_buf[266]*(-4)+in_buf[267]*(-5)+in_buf[268]*(-5)+in_buf[269]*(0)+in_buf[270]*(-3)+in_buf[271]*(-5)+in_buf[272]*(-5)+in_buf[273]*(1)+in_buf[274]*(-2)+in_buf[275]*(-1)+in_buf[276]*(2)+in_buf[277]*(6)+in_buf[278]*(-2)+in_buf[279]*(-1)+in_buf[280]*(2)+in_buf[281]*(4)+in_buf[282]*(2)+in_buf[283]*(1)+in_buf[284]*(-1)+in_buf[285]*(-6)+in_buf[286]*(-3)+in_buf[287]*(-6)+in_buf[288]*(0)+in_buf[289]*(0)+in_buf[290]*(0)+in_buf[291]*(0)+in_buf[292]*(0)+in_buf[293]*(-5)+in_buf[294]*(-2)+in_buf[295]*(3)+in_buf[296]*(-2)+in_buf[297]*(-3)+in_buf[298]*(-5)+in_buf[299]*(1)+in_buf[300]*(0)+in_buf[301]*(-5)+in_buf[302]*(-1)+in_buf[303]*(1)+in_buf[304]*(-4)+in_buf[305]*(-2)+in_buf[306]*(3)+in_buf[307]*(-2)+in_buf[308]*(1)+in_buf[309]*(-1)+in_buf[310]*(0)+in_buf[311]*(3)+in_buf[312]*(-3)+in_buf[313]*(0)+in_buf[314]*(-5)+in_buf[315]*(-2)+in_buf[316]*(0)+in_buf[317]*(-8)+in_buf[318]*(-5)+in_buf[319]*(0)+in_buf[320]*(-1)+in_buf[321]*(-7)+in_buf[322]*(-6)+in_buf[323]*(-1)+in_buf[324]*(-1)+in_buf[325]*(0)+in_buf[326]*(-2)+in_buf[327]*(-1)+in_buf[328]*(-5)+in_buf[329]*(-1)+in_buf[330]*(3)+in_buf[331]*(-1)+in_buf[332]*(0)+in_buf[333]*(3)+in_buf[334]*(-3)+in_buf[335]*(3)+in_buf[336]*(1)+in_buf[337]*(-3)+in_buf[338]*(0)+in_buf[339]*(0)+in_buf[340]*(0)+in_buf[341]*(0)+in_buf[342]*(0)+in_buf[343]*(-6)+in_buf[344]*(-2)+in_buf[345]*(-6)+in_buf[346]*(-2)+in_buf[347]*(0)+in_buf[348]*(-4)+in_buf[349]*(-5)+in_buf[350]*(-6)+in_buf[351]*(2)+in_buf[352]*(-2)+in_buf[353]*(-2)+in_buf[354]*(0)+in_buf[355]*(-2)+in_buf[356]*(-3)+in_buf[357]*(-2)+in_buf[358]*(-1)+in_buf[359]*(0)+in_buf[360]*(-4)+in_buf[361]*(-1)+in_buf[362]*(4)+in_buf[363]*(0)+in_buf[364]*(0)+in_buf[365]*(4)+in_buf[366]*(-1)+in_buf[367]*(-2)+in_buf[368]*(-1)+in_buf[369]*(-3)+in_buf[370]*(0)+in_buf[371]*(-4)+in_buf[372]*(1)+in_buf[373]*(1)+in_buf[374]*(-1)+in_buf[375]*(-3)+in_buf[376]*(-6)+in_buf[377]*(0)+in_buf[378]*(-3)+in_buf[379]*(0)+in_buf[380]*(-5)+in_buf[381]*(-6)+in_buf[382]*(-5)+in_buf[383]*(0)+in_buf[384]*(-5)+in_buf[385]*(-5)+in_buf[386]*(2)+in_buf[387]*(-3)+in_buf[388]*(-3)+in_buf[389]*(2)+in_buf[390]*(1)+in_buf[391]*(0)+in_buf[392]*(-1)+in_buf[393]*(5)+in_buf[394]*(4)+in_buf[395]*(3)+in_buf[396]*(0)+in_buf[397]*(-2)+in_buf[398]*(4)+in_buf[399]*(2)+in_buf[400]*(3)+in_buf[401]*(0)+in_buf[402]*(-2)+in_buf[403]*(0)+in_buf[404]*(2)+in_buf[405]*(1)+in_buf[406]*(-3)+in_buf[407]*(-6)+in_buf[408]*(-5)+in_buf[409]*(0)+in_buf[410]*(-3)+in_buf[411]*(-3)+in_buf[412]*(-5)+in_buf[413]*(-2)+in_buf[414]*(2)+in_buf[415]*(3)+in_buf[416]*(1)+in_buf[417]*(0)+in_buf[418]*(1)+in_buf[419]*(-1)+in_buf[420]*(3)+in_buf[421]*(4)+in_buf[422]*(0)+in_buf[423]*(0)+in_buf[424]*(0)+in_buf[425]*(2)+in_buf[426]*(-1)+in_buf[427]*(-2)+in_buf[428]*(-4)+in_buf[429]*(0)+in_buf[430]*(-1)+in_buf[431]*(0)+in_buf[432]*(-3)+in_buf[433]*(2)+in_buf[434]*(-3)+in_buf[435]*(-1)+in_buf[436]*(-1)+in_buf[437]*(-1)+in_buf[438]*(-1)+in_buf[439]*(2)+in_buf[440]*(-4)+in_buf[441]*(-1)+in_buf[442]*(2)+in_buf[443]*(-4)+in_buf[444]*(0)+in_buf[445]*(3)+in_buf[446]*(0)+in_buf[447]*(1)+in_buf[448]*(-2)+in_buf[449]*(-2)+in_buf[450]*(0)+in_buf[451]*(0)+in_buf[452]*(0)+in_buf[453]*(-2)+in_buf[454]*(-2)+in_buf[455]*(3)+in_buf[456]*(-1)+in_buf[457]*(-5)+in_buf[458]*(2)+in_buf[459]*(-3)+in_buf[460]*(2)+in_buf[461]*(0)+in_buf[462]*(-4)+in_buf[463]*(2)+in_buf[464]*(-4)+in_buf[465]*(-1)+in_buf[466]*(-2)+in_buf[467]*(2)+in_buf[468]*(-2)+in_buf[469]*(2)+in_buf[470]*(0)+in_buf[471]*(-1)+in_buf[472]*(0)+in_buf[473]*(-2)+in_buf[474]*(5)+in_buf[475]*(4)+in_buf[476]*(0)+in_buf[477]*(3)+in_buf[478]*(4)+in_buf[479]*(0)+in_buf[480]*(0)+in_buf[481]*(0)+in_buf[482]*(0)+in_buf[483]*(-1)+in_buf[484]*(-1)+in_buf[485]*(-2)+in_buf[486]*(-2)+in_buf[487]*(3)+in_buf[488]*(-5)+in_buf[489]*(-2)+in_buf[490]*(-2)+in_buf[491]*(-3)+in_buf[492]*(1)+in_buf[493]*(-5)+in_buf[494]*(0)+in_buf[495]*(-3)+in_buf[496]*(-5)+in_buf[497]*(-4)+in_buf[498]*(0)+in_buf[499]*(0)+in_buf[500]*(5)+in_buf[501]*(0)+in_buf[502]*(4)+in_buf[503]*(-3)+in_buf[504]*(0)+in_buf[505]*(0)+in_buf[506]*(1)+in_buf[507]*(-2)+in_buf[508]*(1)+in_buf[509]*(1)+in_buf[510]*(0)+in_buf[511]*(-2)+in_buf[512]*(-1)+in_buf[513]*(-4)+in_buf[514]*(1)+in_buf[515]*(1)+in_buf[516]*(3)+in_buf[517]*(0)+in_buf[518]*(-2)+in_buf[519]*(-3)+in_buf[520]*(-1)+in_buf[521]*(-3)+in_buf[522]*(-2)+in_buf[523]*(-5)+in_buf[524]*(-5)+in_buf[525]*(-4)+in_buf[526]*(-3)+in_buf[527]*(-3)+in_buf[528]*(-1)+in_buf[529]*(3)+in_buf[530]*(-1)+in_buf[531]*(0)+in_buf[532]*(1)+in_buf[533]*(4)+in_buf[534]*(4)+in_buf[535]*(-6)+in_buf[536]*(0)+in_buf[537]*(2)+in_buf[538]*(1)+in_buf[539]*(3)+in_buf[540]*(-3)+in_buf[541]*(-1)+in_buf[542]*(4)+in_buf[543]*(0)+in_buf[544]*(1)+in_buf[545]*(3)+in_buf[546]*(0)+in_buf[547]*(-1)+in_buf[548]*(-6)+in_buf[549]*(2)+in_buf[550]*(-3)+in_buf[551]*(-4)+in_buf[552]*(-1)+in_buf[553]*(2)+in_buf[554]*(0)+in_buf[555]*(-2)+in_buf[556]*(7)+in_buf[557]*(6)+in_buf[558]*(3)+in_buf[559]*(-2)+in_buf[560]*(3)+in_buf[561]*(-1)+in_buf[562]*(3)+in_buf[563]*(-6)+in_buf[564]*(-1)+in_buf[565]*(-2)+in_buf[566]*(0)+in_buf[567]*(3)+in_buf[568]*(0)+in_buf[569]*(3)+in_buf[570]*(-3)+in_buf[571]*(-2)+in_buf[572]*(2)+in_buf[573]*(-1)+in_buf[574]*(1)+in_buf[575]*(-6)+in_buf[576]*(1)+in_buf[577]*(-3)+in_buf[578]*(-2)+in_buf[579]*(-3)+in_buf[580]*(2)+in_buf[581]*(3)+in_buf[582]*(-1)+in_buf[583]*(8)+in_buf[584]*(0)+in_buf[585]*(5)+in_buf[586]*(3)+in_buf[587]*(0)+in_buf[588]*(0)+in_buf[589]*(-1)+in_buf[590]*(3)+in_buf[591]*(-2)+in_buf[592]*(4)+in_buf[593]*(4)+in_buf[594]*(2)+in_buf[595]*(3)+in_buf[596]*(5)+in_buf[597]*(5)+in_buf[598]*(0)+in_buf[599]*(3)+in_buf[600]*(-1)+in_buf[601]*(0)+in_buf[602]*(-3)+in_buf[603]*(0)+in_buf[604]*(0)+in_buf[605]*(0)+in_buf[606]*(4)+in_buf[607]*(2)+in_buf[608]*(-3)+in_buf[609]*(1)+in_buf[610]*(7)+in_buf[611]*(5)+in_buf[612]*(1)+in_buf[613]*(3)+in_buf[614]*(1)+in_buf[615]*(0)+in_buf[616]*(1)+in_buf[617]*(1)+in_buf[618]*(5)+in_buf[619]*(-4)+in_buf[620]*(1)+in_buf[621]*(2)+in_buf[622]*(2)+in_buf[623]*(-2)+in_buf[624]*(-3)+in_buf[625]*(-2)+in_buf[626]*(0)+in_buf[627]*(-3)+in_buf[628]*(1)+in_buf[629]*(0)+in_buf[630]*(0)+in_buf[631]*(0)+in_buf[632]*(-1)+in_buf[633]*(-5)+in_buf[634]*(2)+in_buf[635]*(-4)+in_buf[636]*(-3)+in_buf[637]*(0)+in_buf[638]*(-1)+in_buf[639]*(-1)+in_buf[640]*(0)+in_buf[641]*(3)+in_buf[642]*(-2)+in_buf[643]*(4)+in_buf[644]*(-2)+in_buf[645]*(-2)+in_buf[646]*(3)+in_buf[647]*(0)+in_buf[648]*(-1)+in_buf[649]*(-1)+in_buf[650]*(-3)+in_buf[651]*(0)+in_buf[652]*(0)+in_buf[653]*(-2)+in_buf[654]*(1)+in_buf[655]*(0)+in_buf[656]*(-5)+in_buf[657]*(-2)+in_buf[658]*(-4)+in_buf[659]*(-2)+in_buf[660]*(-6)+in_buf[661]*(-6)+in_buf[662]*(-3)+in_buf[663]*(-6)+in_buf[664]*(2)+in_buf[665]*(3)+in_buf[666]*(2)+in_buf[667]*(6)+in_buf[668]*(1)+in_buf[669]*(0)+in_buf[670]*(-3)+in_buf[671]*(0)+in_buf[672]*(0)+in_buf[673]*(2)+in_buf[674]*(2)+in_buf[675]*(-5)+in_buf[676]*(1)+in_buf[677]*(2)+in_buf[678]*(1)+in_buf[679]*(2)+in_buf[680]*(-4)+in_buf[681]*(-2)+in_buf[682]*(-3)+in_buf[683]*(1)+in_buf[684]*(-1)+in_buf[685]*(-2)+in_buf[686]*(-5)+in_buf[687]*(-6)+in_buf[688]*(-2)+in_buf[689]*(-3)+in_buf[690]*(-2)+in_buf[691]*(-5)+in_buf[692]*(-5)+in_buf[693]*(2)+in_buf[694]*(-2)+in_buf[695]*(0)+in_buf[696]*(1)+in_buf[697]*(0)+in_buf[698]*(0)+in_buf[699]*(-2)+in_buf[700]*(-3)+in_buf[701]*(4)+in_buf[702]*(-3)+in_buf[703]*(0)+in_buf[704]*(-3)+in_buf[705]*(2)+in_buf[706]*(2)+in_buf[707]*(1)+in_buf[708]*(-1)+in_buf[709]*(3)+in_buf[710]*(3)+in_buf[711]*(0)+in_buf[712]*(0)+in_buf[713]*(-2)+in_buf[714]*(0)+in_buf[715]*(0)+in_buf[716]*(-2)+in_buf[717]*(2)+in_buf[718]*(-3)+in_buf[719]*(2)+in_buf[720]*(-2)+in_buf[721]*(0)+in_buf[722]*(3)+in_buf[723]*(0)+in_buf[724]*(4)+in_buf[725]*(3)+in_buf[726]*(0)+in_buf[727]*(-4)+in_buf[728]*(-1)+in_buf[729]*(2)+in_buf[730]*(-1)+in_buf[731]*(-2)+in_buf[732]*(2)+in_buf[733]*(0)+in_buf[734]*(0)+in_buf[735]*(2)+in_buf[736]*(1)+in_buf[737]*(5)+in_buf[738]*(2)+in_buf[739]*(0)+in_buf[740]*(3)+in_buf[741]*(-2)+in_buf[742]*(3)+in_buf[743]*(-3)+in_buf[744]*(-2)+in_buf[745]*(4)+in_buf[746]*(-3)+in_buf[747]*(3)+in_buf[748]*(3)+in_buf[749]*(4)+in_buf[750]*(-3)+in_buf[751]*(3)+in_buf[752]*(-3)+in_buf[753]*(3)+in_buf[754]*(2)+in_buf[755]*(0)+in_buf[756]*(2)+in_buf[757]*(3)+in_buf[758]*(-3)+in_buf[759]*(3)+in_buf[760]*(3)+in_buf[761]*(3)+in_buf[762]*(-2)+in_buf[763]*(2)+in_buf[764]*(3)+in_buf[765]*(1)+in_buf[766]*(3)+in_buf[767]*(5)+in_buf[768]*(-3)+in_buf[769]*(4)+in_buf[770]*(0)+in_buf[771]*(-2)+in_buf[772]*(2)+in_buf[773]*(-2)+in_buf[774]*(1)+in_buf[775]*(0)+in_buf[776]*(2)+in_buf[777]*(2)+in_buf[778]*(4)+in_buf[779]*(3)+in_buf[780]*(0)+in_buf[781]*(0)+in_buf[782]*(0)+in_buf[783]*(4);
assign in_buf_weight010=in_buf[0]*(2)+in_buf[1]*(0)+in_buf[2]*(3)+in_buf[3]*(1)+in_buf[4]*(-2)+in_buf[5]*(0)+in_buf[6]*(3)+in_buf[7]*(3)+in_buf[8]*(0)+in_buf[9]*(0)+in_buf[10]*(-1)+in_buf[11]*(1)+in_buf[12]*(-3)+in_buf[13]*(-4)+in_buf[14]*(0)+in_buf[15]*(6)+in_buf[16]*(0)+in_buf[17]*(-3)+in_buf[18]*(-3)+in_buf[19]*(3)+in_buf[20]*(0)+in_buf[21]*(-1)+in_buf[22]*(2)+in_buf[23]*(0)+in_buf[24]*(-2)+in_buf[25]*(-1)+in_buf[26]*(1)+in_buf[27]*(-3)+in_buf[28]*(-2)+in_buf[29]*(2)+in_buf[30]*(-3)+in_buf[31]*(-2)+in_buf[32]*(1)+in_buf[33]*(-8)+in_buf[34]*(-4)+in_buf[35]*(-5)+in_buf[36]*(-11)+in_buf[37]*(-11)+in_buf[38]*(-7)+in_buf[39]*(-8)+in_buf[40]*(-18)+in_buf[41]*(-4)+in_buf[42]*(16)+in_buf[43]*(-6)+in_buf[44]*(-5)+in_buf[45]*(-13)+in_buf[46]*(-24)+in_buf[47]*(-24)+in_buf[48]*(-18)+in_buf[49]*(-19)+in_buf[50]*(-14)+in_buf[51]*(-13)+in_buf[52]*(0)+in_buf[53]*(0)+in_buf[54]*(-1)+in_buf[55]*(4)+in_buf[56]*(0)+in_buf[57]*(-3)+in_buf[58]*(-1)+in_buf[59]*(-2)+in_buf[60]*(-5)+in_buf[61]*(-3)+in_buf[62]*(-15)+in_buf[63]*(-13)+in_buf[64]*(-17)+in_buf[65]*(-20)+in_buf[66]*(-9)+in_buf[67]*(-31)+in_buf[68]*(-48)+in_buf[69]*(-50)+in_buf[70]*(-42)+in_buf[71]*(-17)+in_buf[72]*(-11)+in_buf[73]*(3)+in_buf[74]*(0)+in_buf[75]*(-13)+in_buf[76]*(-6)+in_buf[77]*(-13)+in_buf[78]*(-21)+in_buf[79]*(-14)+in_buf[80]*(11)+in_buf[81]*(0)+in_buf[82]*(2)+in_buf[83]*(0)+in_buf[84]*(-2)+in_buf[85]*(0)+in_buf[86]*(6)+in_buf[87]*(-11)+in_buf[88]*(-7)+in_buf[89]*(-15)+in_buf[90]*(-26)+in_buf[91]*(-18)+in_buf[92]*(-19)+in_buf[93]*(-20)+in_buf[94]*(-19)+in_buf[95]*(-41)+in_buf[96]*(-59)+in_buf[97]*(-64)+in_buf[98]*(-40)+in_buf[99]*(-20)+in_buf[100]*(-27)+in_buf[101]*(-32)+in_buf[102]*(-5)+in_buf[103]*(-18)+in_buf[104]*(-47)+in_buf[105]*(-30)+in_buf[106]*(-29)+in_buf[107]*(-33)+in_buf[108]*(-27)+in_buf[109]*(-23)+in_buf[110]*(-21)+in_buf[111]*(1)+in_buf[112]*(3)+in_buf[113]*(1)+in_buf[114]*(23)+in_buf[115]*(28)+in_buf[116]*(4)+in_buf[117]*(-9)+in_buf[118]*(-15)+in_buf[119]*(-5)+in_buf[120]*(-9)+in_buf[121]*(-12)+in_buf[122]*(-9)+in_buf[123]*(-11)+in_buf[124]*(-13)+in_buf[125]*(-17)+in_buf[126]*(-12)+in_buf[127]*(-23)+in_buf[128]*(-23)+in_buf[129]*(-14)+in_buf[130]*(6)+in_buf[131]*(-5)+in_buf[132]*(-18)+in_buf[133]*(-32)+in_buf[134]*(-28)+in_buf[135]*(-17)+in_buf[136]*(-12)+in_buf[137]*(-12)+in_buf[138]*(13)+in_buf[139]*(-2)+in_buf[140]*(1)+in_buf[141]*(2)+in_buf[142]*(-10)+in_buf[143]*(-5)+in_buf[144]*(1)+in_buf[145]*(15)+in_buf[146]*(3)+in_buf[147]*(4)+in_buf[148]*(-3)+in_buf[149]*(-8)+in_buf[150]*(-16)+in_buf[151]*(17)+in_buf[152]*(29)+in_buf[153]*(12)+in_buf[154]*(6)+in_buf[155]*(-13)+in_buf[156]*(-15)+in_buf[157]*(3)+in_buf[158]*(-11)+in_buf[159]*(-21)+in_buf[160]*(-19)+in_buf[161]*(-21)+in_buf[162]*(-14)+in_buf[163]*(-15)+in_buf[164]*(-25)+in_buf[165]*(-18)+in_buf[166]*(-21)+in_buf[167]*(-2)+in_buf[168]*(2)+in_buf[169]*(15)+in_buf[170]*(3)+in_buf[171]*(17)+in_buf[172]*(15)+in_buf[173]*(6)+in_buf[174]*(13)+in_buf[175]*(1)+in_buf[176]*(5)+in_buf[177]*(13)+in_buf[178]*(24)+in_buf[179]*(34)+in_buf[180]*(42)+in_buf[181]*(31)+in_buf[182]*(17)+in_buf[183]*(19)+in_buf[184]*(19)+in_buf[185]*(20)+in_buf[186]*(7)+in_buf[187]*(0)+in_buf[188]*(6)+in_buf[189]*(0)+in_buf[190]*(4)+in_buf[191]*(16)+in_buf[192]*(-12)+in_buf[193]*(-4)+in_buf[194]*(-7)+in_buf[195]*(-20)+in_buf[196]*(1)+in_buf[197]*(21)+in_buf[198]*(15)+in_buf[199]*(31)+in_buf[200]*(7)+in_buf[201]*(-23)+in_buf[202]*(1)+in_buf[203]*(-9)+in_buf[204]*(7)+in_buf[205]*(23)+in_buf[206]*(25)+in_buf[207]*(29)+in_buf[208]*(35)+in_buf[209]*(38)+in_buf[210]*(20)+in_buf[211]*(13)+in_buf[212]*(4)+in_buf[213]*(5)+in_buf[214]*(9)+in_buf[215]*(9)+in_buf[216]*(14)+in_buf[217]*(4)+in_buf[218]*(0)+in_buf[219]*(17)+in_buf[220]*(16)+in_buf[221]*(16)+in_buf[222]*(-15)+in_buf[223]*(-26)+in_buf[224]*(-3)+in_buf[225]*(6)+in_buf[226]*(31)+in_buf[227]*(37)+in_buf[228]*(1)+in_buf[229]*(7)+in_buf[230]*(-4)+in_buf[231]*(0)+in_buf[232]*(32)+in_buf[233]*(32)+in_buf[234]*(20)+in_buf[235]*(30)+in_buf[236]*(29)+in_buf[237]*(34)+in_buf[238]*(21)+in_buf[239]*(1)+in_buf[240]*(-9)+in_buf[241]*(-2)+in_buf[242]*(12)+in_buf[243]*(2)+in_buf[244]*(2)+in_buf[245]*(3)+in_buf[246]*(19)+in_buf[247]*(24)+in_buf[248]*(27)+in_buf[249]*(37)+in_buf[250]*(20)+in_buf[251]*(12)+in_buf[252]*(-6)+in_buf[253]*(5)+in_buf[254]*(29)+in_buf[255]*(31)+in_buf[256]*(4)+in_buf[257]*(7)+in_buf[258]*(8)+in_buf[259]*(13)+in_buf[260]*(21)+in_buf[261]*(18)+in_buf[262]*(1)+in_buf[263]*(8)+in_buf[264]*(19)+in_buf[265]*(10)+in_buf[266]*(3)+in_buf[267]*(-19)+in_buf[268]*(-18)+in_buf[269]*(0)+in_buf[270]*(-6)+in_buf[271]*(-9)+in_buf[272]*(8)+in_buf[273]*(10)+in_buf[274]*(25)+in_buf[275]*(32)+in_buf[276]*(9)+in_buf[277]*(10)+in_buf[278]*(41)+in_buf[279]*(33)+in_buf[280]*(-4)+in_buf[281]*(-6)+in_buf[282]*(26)+in_buf[283]*(12)+in_buf[284]*(20)+in_buf[285]*(-10)+in_buf[286]*(9)+in_buf[287]*(5)+in_buf[288]*(-3)+in_buf[289]*(-7)+in_buf[290]*(-18)+in_buf[291]*(-11)+in_buf[292]*(-10)+in_buf[293]*(-16)+in_buf[294]*(-15)+in_buf[295]*(-27)+in_buf[296]*(-18)+in_buf[297]*(-19)+in_buf[298]*(-1)+in_buf[299]*(-7)+in_buf[300]*(7)+in_buf[301]*(1)+in_buf[302]*(26)+in_buf[303]*(36)+in_buf[304]*(9)+in_buf[305]*(14)+in_buf[306]*(3)+in_buf[307]*(30)+in_buf[308]*(5)+in_buf[309]*(-38)+in_buf[310]*(18)+in_buf[311]*(31)+in_buf[312]*(7)+in_buf[313]*(8)+in_buf[314]*(0)+in_buf[315]*(4)+in_buf[316]*(-4)+in_buf[317]*(-15)+in_buf[318]*(-22)+in_buf[319]*(-24)+in_buf[320]*(-10)+in_buf[321]*(-18)+in_buf[322]*(-10)+in_buf[323]*(-5)+in_buf[324]*(11)+in_buf[325]*(-4)+in_buf[326]*(-7)+in_buf[327]*(0)+in_buf[328]*(3)+in_buf[329]*(-4)+in_buf[330]*(4)+in_buf[331]*(6)+in_buf[332]*(12)+in_buf[333]*(23)+in_buf[334]*(8)+in_buf[335]*(3)+in_buf[336]*(11)+in_buf[337]*(-3)+in_buf[338]*(29)+in_buf[339]*(9)+in_buf[340]*(-4)+in_buf[341]*(4)+in_buf[342]*(-14)+in_buf[343]*(-16)+in_buf[344]*(-26)+in_buf[345]*(-37)+in_buf[346]*(-33)+in_buf[347]*(-39)+in_buf[348]*(-22)+in_buf[349]*(6)+in_buf[350]*(10)+in_buf[351]*(16)+in_buf[352]*(8)+in_buf[353]*(5)+in_buf[354]*(17)+in_buf[355]*(11)+in_buf[356]*(6)+in_buf[357]*(6)+in_buf[358]*(1)+in_buf[359]*(9)+in_buf[360]*(-6)+in_buf[361]*(24)+in_buf[362]*(11)+in_buf[363]*(18)+in_buf[364]*(-22)+in_buf[365]*(0)+in_buf[366]*(14)+in_buf[367]*(-7)+in_buf[368]*(0)+in_buf[369]*(-29)+in_buf[370]*(-32)+in_buf[371]*(-32)+in_buf[372]*(-26)+in_buf[373]*(-27)+in_buf[374]*(-19)+in_buf[375]*(-6)+in_buf[376]*(6)+in_buf[377]*(24)+in_buf[378]*(26)+in_buf[379]*(18)+in_buf[380]*(7)+in_buf[381]*(5)+in_buf[382]*(10)+in_buf[383]*(13)+in_buf[384]*(14)+in_buf[385]*(7)+in_buf[386]*(16)+in_buf[387]*(-6)+in_buf[388]*(-20)+in_buf[389]*(19)+in_buf[390]*(11)+in_buf[391]*(24)+in_buf[392]*(-17)+in_buf[393]*(1)+in_buf[394]*(-15)+in_buf[395]*(-15)+in_buf[396]*(7)+in_buf[397]*(-36)+in_buf[398]*(-30)+in_buf[399]*(-22)+in_buf[400]*(-20)+in_buf[401]*(-9)+in_buf[402]*(8)+in_buf[403]*(13)+in_buf[404]*(29)+in_buf[405]*(30)+in_buf[406]*(20)+in_buf[407]*(19)+in_buf[408]*(4)+in_buf[409]*(26)+in_buf[410]*(18)+in_buf[411]*(12)+in_buf[412]*(13)+in_buf[413]*(-2)+in_buf[414]*(2)+in_buf[415]*(-22)+in_buf[416]*(-39)+in_buf[417]*(-17)+in_buf[418]*(-3)+in_buf[419]*(15)+in_buf[420]*(-9)+in_buf[421]*(12)+in_buf[422]*(-13)+in_buf[423]*(-29)+in_buf[424]*(-3)+in_buf[425]*(0)+in_buf[426]*(-28)+in_buf[427]*(-20)+in_buf[428]*(-5)+in_buf[429]*(-2)+in_buf[430]*(16)+in_buf[431]*(19)+in_buf[432]*(18)+in_buf[433]*(23)+in_buf[434]*(26)+in_buf[435]*(33)+in_buf[436]*(14)+in_buf[437]*(36)+in_buf[438]*(15)+in_buf[439]*(3)+in_buf[440]*(7)+in_buf[441]*(-1)+in_buf[442]*(13)+in_buf[443]*(9)+in_buf[444]*(-15)+in_buf[445]*(-40)+in_buf[446]*(36)+in_buf[447]*(6)+in_buf[448]*(6)+in_buf[449]*(22)+in_buf[450]*(24)+in_buf[451]*(-16)+in_buf[452]*(6)+in_buf[453]*(-12)+in_buf[454]*(-4)+in_buf[455]*(6)+in_buf[456]*(11)+in_buf[457]*(14)+in_buf[458]*(9)+in_buf[459]*(2)+in_buf[460]*(20)+in_buf[461]*(33)+in_buf[462]*(28)+in_buf[463]*(16)+in_buf[464]*(17)+in_buf[465]*(25)+in_buf[466]*(10)+in_buf[467]*(-13)+in_buf[468]*(7)+in_buf[469]*(-1)+in_buf[470]*(-6)+in_buf[471]*(0)+in_buf[472]*(-8)+in_buf[473]*(-33)+in_buf[474]*(2)+in_buf[475]*(5)+in_buf[476]*(-2)+in_buf[477]*(15)+in_buf[478]*(19)+in_buf[479]*(-2)+in_buf[480]*(-4)+in_buf[481]*(-13)+in_buf[482]*(-3)+in_buf[483]*(9)+in_buf[484]*(14)+in_buf[485]*(8)+in_buf[486]*(-6)+in_buf[487]*(-1)+in_buf[488]*(8)+in_buf[489]*(24)+in_buf[490]*(13)+in_buf[491]*(6)+in_buf[492]*(3)+in_buf[493]*(3)+in_buf[494]*(-9)+in_buf[495]*(-19)+in_buf[496]*(-9)+in_buf[497]*(-6)+in_buf[498]*(-21)+in_buf[499]*(-11)+in_buf[500]*(-3)+in_buf[501]*(0)+in_buf[502]*(16)+in_buf[503]*(-12)+in_buf[504]*(17)+in_buf[505]*(10)+in_buf[506]*(26)+in_buf[507]*(-6)+in_buf[508]*(-18)+in_buf[509]*(-4)+in_buf[510]*(8)+in_buf[511]*(-8)+in_buf[512]*(-5)+in_buf[513]*(-12)+in_buf[514]*(-8)+in_buf[515]*(-11)+in_buf[516]*(-22)+in_buf[517]*(0)+in_buf[518]*(-4)+in_buf[519]*(-11)+in_buf[520]*(-9)+in_buf[521]*(-8)+in_buf[522]*(-16)+in_buf[523]*(-14)+in_buf[524]*(-8)+in_buf[525]*(-18)+in_buf[526]*(-17)+in_buf[527]*(-8)+in_buf[528]*(-14)+in_buf[529]*(-6)+in_buf[530]*(33)+in_buf[531]*(-5)+in_buf[532]*(-19)+in_buf[533]*(-32)+in_buf[534]*(23)+in_buf[535]*(-18)+in_buf[536]*(-1)+in_buf[537]*(-8)+in_buf[538]*(-7)+in_buf[539]*(7)+in_buf[540]*(-21)+in_buf[541]*(-17)+in_buf[542]*(-24)+in_buf[543]*(-37)+in_buf[544]*(-36)+in_buf[545]*(-19)+in_buf[546]*(-12)+in_buf[547]*(-15)+in_buf[548]*(-2)+in_buf[549]*(-5)+in_buf[550]*(-12)+in_buf[551]*(-4)+in_buf[552]*(-22)+in_buf[553]*(-22)+in_buf[554]*(-14)+in_buf[555]*(-4)+in_buf[556]*(-33)+in_buf[557]*(-37)+in_buf[558]*(-6)+in_buf[559]*(-16)+in_buf[560]*(4)+in_buf[561]*(-14)+in_buf[562]*(7)+in_buf[563]*(-16)+in_buf[564]*(4)+in_buf[565]*(0)+in_buf[566]*(0)+in_buf[567]*(2)+in_buf[568]*(-6)+in_buf[569]*(-2)+in_buf[570]*(-8)+in_buf[571]*(-26)+in_buf[572]*(-32)+in_buf[573]*(-13)+in_buf[574]*(-12)+in_buf[575]*(-12)+in_buf[576]*(2)+in_buf[577]*(-18)+in_buf[578]*(-14)+in_buf[579]*(0)+in_buf[580]*(-19)+in_buf[581]*(-12)+in_buf[582]*(-1)+in_buf[583]*(5)+in_buf[584]*(-15)+in_buf[585]*(-32)+in_buf[586]*(-20)+in_buf[587]*(-5)+in_buf[588]*(-14)+in_buf[589]*(20)+in_buf[590]*(18)+in_buf[591]*(-13)+in_buf[592]*(3)+in_buf[593]*(0)+in_buf[594]*(-2)+in_buf[595]*(6)+in_buf[596]*(12)+in_buf[597]*(-2)+in_buf[598]*(0)+in_buf[599]*(-3)+in_buf[600]*(-10)+in_buf[601]*(-7)+in_buf[602]*(-8)+in_buf[603]*(-9)+in_buf[604]*(-8)+in_buf[605]*(-29)+in_buf[606]*(-41)+in_buf[607]*(-29)+in_buf[608]*(-30)+in_buf[609]*(-15)+in_buf[610]*(4)+in_buf[611]*(-5)+in_buf[612]*(-36)+in_buf[613]*(-38)+in_buf[614]*(-35)+in_buf[615]*(-3)+in_buf[616]*(-20)+in_buf[617]*(17)+in_buf[618]*(15)+in_buf[619]*(-22)+in_buf[620]*(25)+in_buf[621]*(11)+in_buf[622]*(11)+in_buf[623]*(18)+in_buf[624]*(17)+in_buf[625]*(-7)+in_buf[626]*(1)+in_buf[627]*(9)+in_buf[628]*(4)+in_buf[629]*(0)+in_buf[630]*(-2)+in_buf[631]*(-11)+in_buf[632]*(-25)+in_buf[633]*(-43)+in_buf[634]*(-42)+in_buf[635]*(-29)+in_buf[636]*(-16)+in_buf[637]*(-15)+in_buf[638]*(17)+in_buf[639]*(-4)+in_buf[640]*(-23)+in_buf[641]*(0)+in_buf[642]*(-27)+in_buf[643]*(-2)+in_buf[644]*(4)+in_buf[645]*(-2)+in_buf[646]*(21)+in_buf[647]*(0)+in_buf[648]*(28)+in_buf[649]*(8)+in_buf[650]*(18)+in_buf[651]*(23)+in_buf[652]*(7)+in_buf[653]*(-11)+in_buf[654]*(-1)+in_buf[655]*(10)+in_buf[656]*(6)+in_buf[657]*(16)+in_buf[658]*(12)+in_buf[659]*(-2)+in_buf[660]*(-20)+in_buf[661]*(-33)+in_buf[662]*(-23)+in_buf[663]*(-22)+in_buf[664]*(3)+in_buf[665]*(-6)+in_buf[666]*(-10)+in_buf[667]*(-11)+in_buf[668]*(-11)+in_buf[669]*(0)+in_buf[670]*(-35)+in_buf[671]*(0)+in_buf[672]*(0)+in_buf[673]*(3)+in_buf[674]*(14)+in_buf[675]*(23)+in_buf[676]*(56)+in_buf[677]*(23)+in_buf[678]*(39)+in_buf[679]*(21)+in_buf[680]*(15)+in_buf[681]*(-8)+in_buf[682]*(5)+in_buf[683]*(13)+in_buf[684]*(0)+in_buf[685]*(22)+in_buf[686]*(12)+in_buf[687]*(3)+in_buf[688]*(-10)+in_buf[689]*(-28)+in_buf[690]*(-28)+in_buf[691]*(-4)+in_buf[692]*(15)+in_buf[693]*(0)+in_buf[694]*(-33)+in_buf[695]*(-8)+in_buf[696]*(-39)+in_buf[697]*(-40)+in_buf[698]*(-21)+in_buf[699]*(3)+in_buf[700]*(3)+in_buf[701]*(0)+in_buf[702]*(-4)+in_buf[703]*(1)+in_buf[704]*(23)+in_buf[705]*(65)+in_buf[706]*(34)+in_buf[707]*(25)+in_buf[708]*(20)+in_buf[709]*(22)+in_buf[710]*(33)+in_buf[711]*(14)+in_buf[712]*(0)+in_buf[713]*(12)+in_buf[714]*(22)+in_buf[715]*(2)+in_buf[716]*(0)+in_buf[717]*(-7)+in_buf[718]*(-3)+in_buf[719]*(7)+in_buf[720]*(4)+in_buf[721]*(-27)+in_buf[722]*(-26)+in_buf[723]*(-9)+in_buf[724]*(-14)+in_buf[725]*(-14)+in_buf[726]*(-13)+in_buf[727]*(-1)+in_buf[728]*(-1)+in_buf[729]*(1)+in_buf[730]*(0)+in_buf[731]*(8)+in_buf[732]*(18)+in_buf[733]*(25)+in_buf[734]*(37)+in_buf[735]*(53)+in_buf[736]*(36)+in_buf[737]*(37)+in_buf[738]*(48)+in_buf[739]*(31)+in_buf[740]*(7)+in_buf[741]*(25)+in_buf[742]*(59)+in_buf[743]*(16)+in_buf[744]*(29)+in_buf[745]*(56)+in_buf[746]*(31)+in_buf[747]*(21)+in_buf[748]*(37)+in_buf[749]*(3)+in_buf[750]*(-6)+in_buf[751]*(-2)+in_buf[752]*(1)+in_buf[753]*(3)+in_buf[754]*(3)+in_buf[755]*(-3)+in_buf[756]*(-2)+in_buf[757]*(2)+in_buf[758]*(2)+in_buf[759]*(2)+in_buf[760]*(-14)+in_buf[761]*(-3)+in_buf[762]*(12)+in_buf[763]*(17)+in_buf[764]*(11)+in_buf[765]*(7)+in_buf[766]*(47)+in_buf[767]*(21)+in_buf[768]*(23)+in_buf[769]*(23)+in_buf[770]*(65)+in_buf[771]*(31)+in_buf[772]*(10)+in_buf[773]*(-4)+in_buf[774]*(-2)+in_buf[775]*(7)+in_buf[776]*(0)+in_buf[777]*(7)+in_buf[778]*(-8)+in_buf[779]*(2)+in_buf[780]*(3)+in_buf[781]*(1)+in_buf[782]*(2)+in_buf[783]*(2);
assign in_buf_weight011=in_buf[0]*(0)+in_buf[1]*(-3)+in_buf[2]*(-2)+in_buf[3]*(1)+in_buf[4]*(3)+in_buf[5]*(1)+in_buf[6]*(2)+in_buf[7]*(4)+in_buf[8]*(3)+in_buf[9]*(-1)+in_buf[10]*(-3)+in_buf[11]*(0)+in_buf[12]*(-9)+in_buf[13]*(-3)+in_buf[14]*(22)+in_buf[15]*(14)+in_buf[16]*(-2)+in_buf[17]*(0)+in_buf[18]*(1)+in_buf[19]*(1)+in_buf[20]*(-3)+in_buf[21]*(-4)+in_buf[22]*(3)+in_buf[23]*(2)+in_buf[24]*(-2)+in_buf[25]*(-3)+in_buf[26]*(-2)+in_buf[27]*(-1)+in_buf[28]*(4)+in_buf[29]*(0)+in_buf[30]*(0)+in_buf[31]*(0)+in_buf[32]*(-3)+in_buf[33]*(4)+in_buf[34]*(6)+in_buf[35]*(7)+in_buf[36]*(7)+in_buf[37]*(11)+in_buf[38]*(10)+in_buf[39]*(10)+in_buf[40]*(12)+in_buf[41]*(-17)+in_buf[42]*(-9)+in_buf[43]*(24)+in_buf[44]*(37)+in_buf[45]*(27)+in_buf[46]*(-8)+in_buf[47]*(2)+in_buf[48]*(2)+in_buf[49]*(-4)+in_buf[50]*(0)+in_buf[51]*(8)+in_buf[52]*(2)+in_buf[53]*(2)+in_buf[54]*(0)+in_buf[55]*(-3)+in_buf[56]*(-2)+in_buf[57]*(2)+in_buf[58]*(0)+in_buf[59]*(28)+in_buf[60]*(24)+in_buf[61]*(9)+in_buf[62]*(6)+in_buf[63]*(6)+in_buf[64]*(29)+in_buf[65]*(57)+in_buf[66]*(60)+in_buf[67]*(46)+in_buf[68]*(29)+in_buf[69]*(8)+in_buf[70]*(17)+in_buf[71]*(17)+in_buf[72]*(15)+in_buf[73]*(5)+in_buf[74]*(17)+in_buf[75]*(-1)+in_buf[76]*(16)+in_buf[77]*(19)+in_buf[78]*(9)+in_buf[79]*(4)+in_buf[80]*(18)+in_buf[81]*(12)+in_buf[82]*(-3)+in_buf[83]*(3)+in_buf[84]*(-1)+in_buf[85]*(3)+in_buf[86]*(-2)+in_buf[87]*(26)+in_buf[88]*(-1)+in_buf[89]*(19)+in_buf[90]*(38)+in_buf[91]*(11)+in_buf[92]*(33)+in_buf[93]*(41)+in_buf[94]*(28)+in_buf[95]*(34)+in_buf[96]*(24)+in_buf[97]*(25)+in_buf[98]*(0)+in_buf[99]*(12)+in_buf[100]*(16)+in_buf[101]*(3)+in_buf[102]*(19)+in_buf[103]*(5)+in_buf[104]*(-26)+in_buf[105]*(2)+in_buf[106]*(16)+in_buf[107]*(23)+in_buf[108]*(1)+in_buf[109]*(-17)+in_buf[110]*(-34)+in_buf[111]*(2)+in_buf[112]*(-2)+in_buf[113]*(2)+in_buf[114]*(8)+in_buf[115]*(-25)+in_buf[116]*(-3)+in_buf[117]*(13)+in_buf[118]*(8)+in_buf[119]*(11)+in_buf[120]*(27)+in_buf[121]*(28)+in_buf[122]*(26)+in_buf[123]*(21)+in_buf[124]*(24)+in_buf[125]*(6)+in_buf[126]*(19)+in_buf[127]*(20)+in_buf[128]*(26)+in_buf[129]*(20)+in_buf[130]*(-10)+in_buf[131]*(-2)+in_buf[132]*(-8)+in_buf[133]*(-28)+in_buf[134]*(-22)+in_buf[135]*(-19)+in_buf[136]*(-10)+in_buf[137]*(-6)+in_buf[138]*(20)+in_buf[139]*(1)+in_buf[140]*(-3)+in_buf[141]*(-3)+in_buf[142]*(52)+in_buf[143]*(3)+in_buf[144]*(9)+in_buf[145]*(-29)+in_buf[146]*(-12)+in_buf[147]*(5)+in_buf[148]*(-8)+in_buf[149]*(-4)+in_buf[150]*(3)+in_buf[151]*(14)+in_buf[152]*(18)+in_buf[153]*(4)+in_buf[154]*(6)+in_buf[155]*(8)+in_buf[156]*(18)+in_buf[157]*(23)+in_buf[158]*(-1)+in_buf[159]*(12)+in_buf[160]*(8)+in_buf[161]*(1)+in_buf[162]*(-5)+in_buf[163]*(-20)+in_buf[164]*(0)+in_buf[165]*(7)+in_buf[166]*(14)+in_buf[167]*(-12)+in_buf[168]*(0)+in_buf[169]*(19)+in_buf[170]*(0)+in_buf[171]*(-32)+in_buf[172]*(-14)+in_buf[173]*(-42)+in_buf[174]*(-25)+in_buf[175]*(-11)+in_buf[176]*(-6)+in_buf[177]*(5)+in_buf[178]*(14)+in_buf[179]*(12)+in_buf[180]*(10)+in_buf[181]*(7)+in_buf[182]*(5)+in_buf[183]*(5)+in_buf[184]*(1)+in_buf[185]*(11)+in_buf[186]*(-2)+in_buf[187]*(2)+in_buf[188]*(-6)+in_buf[189]*(-10)+in_buf[190]*(-16)+in_buf[191]*(-18)+in_buf[192]*(-29)+in_buf[193]*(17)+in_buf[194]*(3)+in_buf[195]*(-22)+in_buf[196]*(-4)+in_buf[197]*(-4)+in_buf[198]*(7)+in_buf[199]*(-36)+in_buf[200]*(9)+in_buf[201]*(-19)+in_buf[202]*(-10)+in_buf[203]*(-4)+in_buf[204]*(16)+in_buf[205]*(7)+in_buf[206]*(13)+in_buf[207]*(0)+in_buf[208]*(-1)+in_buf[209]*(3)+in_buf[210]*(2)+in_buf[211]*(10)+in_buf[212]*(-4)+in_buf[213]*(-3)+in_buf[214]*(4)+in_buf[215]*(8)+in_buf[216]*(-10)+in_buf[217]*(7)+in_buf[218]*(0)+in_buf[219]*(-24)+in_buf[220]*(-18)+in_buf[221]*(5)+in_buf[222]*(-14)+in_buf[223]*(-30)+in_buf[224]*(14)+in_buf[225]*(-26)+in_buf[226]*(4)+in_buf[227]*(12)+in_buf[228]*(27)+in_buf[229]*(-9)+in_buf[230]*(-4)+in_buf[231]*(-2)+in_buf[232]*(2)+in_buf[233]*(-3)+in_buf[234]*(4)+in_buf[235]*(-8)+in_buf[236]*(-8)+in_buf[237]*(4)+in_buf[238]*(5)+in_buf[239]*(0)+in_buf[240]*(4)+in_buf[241]*(-1)+in_buf[242]*(8)+in_buf[243]*(15)+in_buf[244]*(0)+in_buf[245]*(7)+in_buf[246]*(1)+in_buf[247]*(-9)+in_buf[248]*(-26)+in_buf[249]*(-3)+in_buf[250]*(-2)+in_buf[251]*(13)+in_buf[252]*(-8)+in_buf[253]*(-27)+in_buf[254]*(11)+in_buf[255]*(25)+in_buf[256]*(13)+in_buf[257]*(-12)+in_buf[258]*(3)+in_buf[259]*(0)+in_buf[260]*(-2)+in_buf[261]*(5)+in_buf[262]*(-2)+in_buf[263]*(-10)+in_buf[264]*(-7)+in_buf[265]*(0)+in_buf[266]*(0)+in_buf[267]*(-7)+in_buf[268]*(-4)+in_buf[269]*(-4)+in_buf[270]*(-1)+in_buf[271]*(14)+in_buf[272]*(3)+in_buf[273]*(1)+in_buf[274]*(0)+in_buf[275]*(1)+in_buf[276]*(-23)+in_buf[277]*(3)+in_buf[278]*(-4)+in_buf[279]*(-22)+in_buf[280]*(-12)+in_buf[281]*(-21)+in_buf[282]*(-18)+in_buf[283]*(17)+in_buf[284]*(11)+in_buf[285]*(16)+in_buf[286]*(25)+in_buf[287]*(3)+in_buf[288]*(-1)+in_buf[289]*(-6)+in_buf[290]*(-6)+in_buf[291]*(-3)+in_buf[292]*(3)+in_buf[293]*(-9)+in_buf[294]*(-7)+in_buf[295]*(-32)+in_buf[296]*(-26)+in_buf[297]*(-15)+in_buf[298]*(0)+in_buf[299]*(3)+in_buf[300]*(0)+in_buf[301]*(3)+in_buf[302]*(4)+in_buf[303]*(25)+in_buf[304]*(-18)+in_buf[305]*(-40)+in_buf[306]*(-11)+in_buf[307]*(0)+in_buf[308]*(-13)+in_buf[309]*(-30)+in_buf[310]*(-12)+in_buf[311]*(15)+in_buf[312]*(20)+in_buf[313]*(24)+in_buf[314]*(15)+in_buf[315]*(4)+in_buf[316]*(-6)+in_buf[317]*(-1)+in_buf[318]*(-13)+in_buf[319]*(-16)+in_buf[320]*(-6)+in_buf[321]*(-8)+in_buf[322]*(2)+in_buf[323]*(-20)+in_buf[324]*(-19)+in_buf[325]*(-15)+in_buf[326]*(-2)+in_buf[327]*(7)+in_buf[328]*(13)+in_buf[329]*(22)+in_buf[330]*(24)+in_buf[331]*(30)+in_buf[332]*(20)+in_buf[333]*(7)+in_buf[334]*(14)+in_buf[335]*(-30)+in_buf[336]*(-17)+in_buf[337]*(-4)+in_buf[338]*(9)+in_buf[339]*(3)+in_buf[340]*(26)+in_buf[341]*(11)+in_buf[342]*(-2)+in_buf[343]*(-3)+in_buf[344]*(-20)+in_buf[345]*(-4)+in_buf[346]*(-21)+in_buf[347]*(-22)+in_buf[348]*(-18)+in_buf[349]*(-9)+in_buf[350]*(1)+in_buf[351]*(0)+in_buf[352]*(-1)+in_buf[353]*(2)+in_buf[354]*(-8)+in_buf[355]*(14)+in_buf[356]*(19)+in_buf[357]*(25)+in_buf[358]*(16)+in_buf[359]*(28)+in_buf[360]*(39)+in_buf[361]*(11)+in_buf[362]*(0)+in_buf[363]*(-26)+in_buf[364]*(21)+in_buf[365]*(-8)+in_buf[366]*(-15)+in_buf[367]*(0)+in_buf[368]*(-10)+in_buf[369]*(-5)+in_buf[370]*(-18)+in_buf[371]*(-13)+in_buf[372]*(-10)+in_buf[373]*(-3)+in_buf[374]*(-16)+in_buf[375]*(-5)+in_buf[376]*(5)+in_buf[377]*(15)+in_buf[378]*(23)+in_buf[379]*(24)+in_buf[380]*(9)+in_buf[381]*(-4)+in_buf[382]*(-6)+in_buf[383]*(14)+in_buf[384]*(21)+in_buf[385]*(16)+in_buf[386]*(36)+in_buf[387]*(28)+in_buf[388]*(11)+in_buf[389]*(20)+in_buf[390]*(42)+in_buf[391]*(21)+in_buf[392]*(-14)+in_buf[393]*(-12)+in_buf[394]*(-21)+in_buf[395]*(0)+in_buf[396]*(-18)+in_buf[397]*(-21)+in_buf[398]*(-6)+in_buf[399]*(-10)+in_buf[400]*(-11)+in_buf[401]*(-3)+in_buf[402]*(10)+in_buf[403]*(24)+in_buf[404]*(11)+in_buf[405]*(30)+in_buf[406]*(18)+in_buf[407]*(16)+in_buf[408]*(15)+in_buf[409]*(0)+in_buf[410]*(5)+in_buf[411]*(1)+in_buf[412]*(6)+in_buf[413]*(18)+in_buf[414]*(19)+in_buf[415]*(-14)+in_buf[416]*(-6)+in_buf[417]*(19)+in_buf[418]*(47)+in_buf[419]*(17)+in_buf[420]*(-18)+in_buf[421]*(-6)+in_buf[422]*(-1)+in_buf[423]*(15)+in_buf[424]*(-19)+in_buf[425]*(-10)+in_buf[426]*(-3)+in_buf[427]*(-9)+in_buf[428]*(11)+in_buf[429]*(15)+in_buf[430]*(14)+in_buf[431]*(23)+in_buf[432]*(13)+in_buf[433]*(33)+in_buf[434]*(27)+in_buf[435]*(8)+in_buf[436]*(14)+in_buf[437]*(-7)+in_buf[438]*(0)+in_buf[439]*(8)+in_buf[440]*(-1)+in_buf[441]*(-5)+in_buf[442]*(-13)+in_buf[443]*(-23)+in_buf[444]*(5)+in_buf[445]*(5)+in_buf[446]*(-2)+in_buf[447]*(37)+in_buf[448]*(1)+in_buf[449]*(5)+in_buf[450]*(2)+in_buf[451]*(-2)+in_buf[452]*(-14)+in_buf[453]*(-11)+in_buf[454]*(6)+in_buf[455]*(-8)+in_buf[456]*(-3)+in_buf[457]*(17)+in_buf[458]*(24)+in_buf[459]*(17)+in_buf[460]*(20)+in_buf[461]*(18)+in_buf[462]*(19)+in_buf[463]*(6)+in_buf[464]*(4)+in_buf[465]*(-1)+in_buf[466]*(0)+in_buf[467]*(-6)+in_buf[468]*(-19)+in_buf[469]*(-11)+in_buf[470]*(-12)+in_buf[471]*(-18)+in_buf[472]*(-1)+in_buf[473]*(31)+in_buf[474]*(30)+in_buf[475]*(31)+in_buf[476]*(-4)+in_buf[477]*(-4)+in_buf[478]*(-9)+in_buf[479]*(11)+in_buf[480]*(-7)+in_buf[481]*(-16)+in_buf[482]*(-7)+in_buf[483]*(-8)+in_buf[484]*(9)+in_buf[485]*(7)+in_buf[486]*(15)+in_buf[487]*(11)+in_buf[488]*(20)+in_buf[489]*(21)+in_buf[490]*(5)+in_buf[491]*(-7)+in_buf[492]*(-7)+in_buf[493]*(-13)+in_buf[494]*(-14)+in_buf[495]*(-6)+in_buf[496]*(-12)+in_buf[497]*(-12)+in_buf[498]*(-5)+in_buf[499]*(-10)+in_buf[500]*(-1)+in_buf[501]*(25)+in_buf[502]*(20)+in_buf[503]*(44)+in_buf[504]*(30)+in_buf[505]*(-7)+in_buf[506]*(0)+in_buf[507]*(7)+in_buf[508]*(0)+in_buf[509]*(-6)+in_buf[510]*(0)+in_buf[511]*(10)+in_buf[512]*(6)+in_buf[513]*(4)+in_buf[514]*(11)+in_buf[515]*(1)+in_buf[516]*(5)+in_buf[517]*(4)+in_buf[518]*(5)+in_buf[519]*(-8)+in_buf[520]*(-7)+in_buf[521]*(-7)+in_buf[522]*(-9)+in_buf[523]*(-2)+in_buf[524]*(2)+in_buf[525]*(-5)+in_buf[526]*(-1)+in_buf[527]*(12)+in_buf[528]*(18)+in_buf[529]*(49)+in_buf[530]*(12)+in_buf[531]*(25)+in_buf[532]*(11)+in_buf[533]*(-24)+in_buf[534]*(-13)+in_buf[535]*(-13)+in_buf[536]*(9)+in_buf[537]*(9)+in_buf[538]*(-6)+in_buf[539]*(8)+in_buf[540]*(5)+in_buf[541]*(2)+in_buf[542]*(16)+in_buf[543]*(-10)+in_buf[544]*(-13)+in_buf[545]*(-1)+in_buf[546]*(-10)+in_buf[547]*(-6)+in_buf[548]*(4)+in_buf[549]*(8)+in_buf[550]*(5)+in_buf[551]*(12)+in_buf[552]*(6)+in_buf[553]*(-6)+in_buf[554]*(28)+in_buf[555]*(38)+in_buf[556]*(8)+in_buf[557]*(58)+in_buf[558]*(56)+in_buf[559]*(16)+in_buf[560]*(0)+in_buf[561]*(-19)+in_buf[562]*(4)+in_buf[563]*(9)+in_buf[564]*(18)+in_buf[565]*(19)+in_buf[566]*(8)+in_buf[567]*(19)+in_buf[568]*(1)+in_buf[569]*(0)+in_buf[570]*(17)+in_buf[571]*(5)+in_buf[572]*(-8)+in_buf[573]*(-5)+in_buf[574]*(0)+in_buf[575]*(6)+in_buf[576]*(1)+in_buf[577]*(0)+in_buf[578]*(18)+in_buf[579]*(3)+in_buf[580]*(17)+in_buf[581]*(11)+in_buf[582]*(16)+in_buf[583]*(21)+in_buf[584]*(2)+in_buf[585]*(40)+in_buf[586]*(45)+in_buf[587]*(6)+in_buf[588]*(-10)+in_buf[589]*(9)+in_buf[590]*(34)+in_buf[591]*(38)+in_buf[592]*(24)+in_buf[593]*(10)+in_buf[594]*(20)+in_buf[595]*(22)+in_buf[596]*(0)+in_buf[597]*(10)+in_buf[598]*(5)+in_buf[599]*(6)+in_buf[600]*(-1)+in_buf[601]*(6)+in_buf[602]*(8)+in_buf[603]*(0)+in_buf[604]*(0)+in_buf[605]*(10)+in_buf[606]*(10)+in_buf[607]*(11)+in_buf[608]*(0)+in_buf[609]*(0)+in_buf[610]*(15)+in_buf[611]*(20)+in_buf[612]*(-12)+in_buf[613]*(18)+in_buf[614]*(10)+in_buf[615]*(-1)+in_buf[616]*(-10)+in_buf[617]*(0)+in_buf[618]*(33)+in_buf[619]*(19)+in_buf[620]*(32)+in_buf[621]*(16)+in_buf[622]*(18)+in_buf[623]*(18)+in_buf[624]*(11)+in_buf[625]*(7)+in_buf[626]*(2)+in_buf[627]*(12)+in_buf[628]*(12)+in_buf[629]*(18)+in_buf[630]*(12)+in_buf[631]*(-8)+in_buf[632]*(-4)+in_buf[633]*(10)+in_buf[634]*(1)+in_buf[635]*(-5)+in_buf[636]*(10)+in_buf[637]*(-4)+in_buf[638]*(1)+in_buf[639]*(10)+in_buf[640]*(9)+in_buf[641]*(17)+in_buf[642]*(-21)+in_buf[643]*(-4)+in_buf[644]*(3)+in_buf[645]*(0)+in_buf[646]*(27)+in_buf[647]*(2)+in_buf[648]*(9)+in_buf[649]*(-3)+in_buf[650]*(-9)+in_buf[651]*(-3)+in_buf[652]*(11)+in_buf[653]*(2)+in_buf[654]*(-10)+in_buf[655]*(1)+in_buf[656]*(10)+in_buf[657]*(25)+in_buf[658]*(0)+in_buf[659]*(3)+in_buf[660]*(0)+in_buf[661]*(5)+in_buf[662]*(16)+in_buf[663]*(1)+in_buf[664]*(12)+in_buf[665]*(16)+in_buf[666]*(40)+in_buf[667]*(34)+in_buf[668]*(10)+in_buf[669]*(12)+in_buf[670]*(-24)+in_buf[671]*(-3)+in_buf[672]*(-3)+in_buf[673]*(0)+in_buf[674]*(-4)+in_buf[675]*(-21)+in_buf[676]*(-13)+in_buf[677]*(-20)+in_buf[678]*(-5)+in_buf[679]*(-9)+in_buf[680]*(1)+in_buf[681]*(-2)+in_buf[682]*(7)+in_buf[683]*(4)+in_buf[684]*(23)+in_buf[685]*(15)+in_buf[686]*(6)+in_buf[687]*(-4)+in_buf[688]*(-2)+in_buf[689]*(-15)+in_buf[690]*(0)+in_buf[691]*(13)+in_buf[692]*(21)+in_buf[693]*(11)+in_buf[694]*(11)+in_buf[695]*(13)+in_buf[696]*(27)+in_buf[697]*(6)+in_buf[698]*(1)+in_buf[699]*(-2)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(10)+in_buf[703]*(-23)+in_buf[704]*(-42)+in_buf[705]*(-35)+in_buf[706]*(1)+in_buf[707]*(18)+in_buf[708]*(12)+in_buf[709]*(10)+in_buf[710]*(8)+in_buf[711]*(-3)+in_buf[712]*(7)+in_buf[713]*(11)+in_buf[714]*(21)+in_buf[715]*(-4)+in_buf[716]*(-1)+in_buf[717]*(17)+in_buf[718]*(17)+in_buf[719]*(21)+in_buf[720]*(21)+in_buf[721]*(7)+in_buf[722]*(-15)+in_buf[723]*(-18)+in_buf[724]*(-4)+in_buf[725]*(3)+in_buf[726]*(5)+in_buf[727]*(2)+in_buf[728]*(1)+in_buf[729]*(4)+in_buf[730]*(1)+in_buf[731]*(3)+in_buf[732]*(25)+in_buf[733]*(6)+in_buf[734]*(3)+in_buf[735]*(23)+in_buf[736]*(23)+in_buf[737]*(7)+in_buf[738]*(-2)+in_buf[739]*(0)+in_buf[740]*(20)+in_buf[741]*(27)+in_buf[742]*(27)+in_buf[743]*(-18)+in_buf[744]*(13)+in_buf[745]*(27)+in_buf[746]*(35)+in_buf[747]*(22)+in_buf[748]*(10)+in_buf[749]*(-2)+in_buf[750]*(12)+in_buf[751]*(21)+in_buf[752]*(24)+in_buf[753]*(-13)+in_buf[754]*(0)+in_buf[755]*(0)+in_buf[756]*(-2)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(0)+in_buf[760]*(-28)+in_buf[761]*(-13)+in_buf[762]*(6)+in_buf[763]*(13)+in_buf[764]*(-1)+in_buf[765]*(13)+in_buf[766]*(-2)+in_buf[767]*(23)+in_buf[768]*(23)+in_buf[769]*(5)+in_buf[770]*(36)+in_buf[771]*(6)+in_buf[772]*(-8)+in_buf[773]*(-11)+in_buf[774]*(-10)+in_buf[775]*(18)+in_buf[776]*(4)+in_buf[777]*(-4)+in_buf[778]*(-11)+in_buf[779]*(-9)+in_buf[780]*(-3)+in_buf[781]*(-3)+in_buf[782]*(4)+in_buf[783]*(-2);
assign in_buf_weight012=in_buf[0]*(-2)+in_buf[1]*(-1)+in_buf[2]*(4)+in_buf[3]*(3)+in_buf[4]*(-2)+in_buf[5]*(4)+in_buf[6]*(-1)+in_buf[7]*(1)+in_buf[8]*(0)+in_buf[9]*(1)+in_buf[10]*(0)+in_buf[11]*(-1)+in_buf[12]*(-2)+in_buf[13]*(2)+in_buf[14]*(-2)+in_buf[15]*(4)+in_buf[16]*(2)+in_buf[17]*(3)+in_buf[18]*(0)+in_buf[19]*(3)+in_buf[20]*(2)+in_buf[21]*(2)+in_buf[22]*(0)+in_buf[23]*(2)+in_buf[24]*(2)+in_buf[25]*(0)+in_buf[26]*(2)+in_buf[27]*(0)+in_buf[28]*(1)+in_buf[29]*(2)+in_buf[30]*(-3)+in_buf[31]*(0)+in_buf[32]*(-3)+in_buf[33]*(-3)+in_buf[34]*(-6)+in_buf[35]*(0)+in_buf[36]*(-1)+in_buf[37]*(-6)+in_buf[38]*(-8)+in_buf[39]*(-2)+in_buf[40]*(-9)+in_buf[41]*(-15)+in_buf[42]*(-1)+in_buf[43]*(5)+in_buf[44]*(0)+in_buf[45]*(-1)+in_buf[46]*(-5)+in_buf[47]*(-6)+in_buf[48]*(1)+in_buf[49]*(2)+in_buf[50]*(1)+in_buf[51]*(-1)+in_buf[52]*(-1)+in_buf[53]*(2)+in_buf[54]*(-1)+in_buf[55]*(0)+in_buf[56]*(0)+in_buf[57]*(-2)+in_buf[58]*(-1)+in_buf[59]*(-12)+in_buf[60]*(-6)+in_buf[61]*(-4)+in_buf[62]*(-3)+in_buf[63]*(-19)+in_buf[64]*(-1)+in_buf[65]*(2)+in_buf[66]*(11)+in_buf[67]*(-18)+in_buf[68]*(-7)+in_buf[69]*(-35)+in_buf[70]*(-26)+in_buf[71]*(-16)+in_buf[72]*(-20)+in_buf[73]*(-5)+in_buf[74]*(14)+in_buf[75]*(14)+in_buf[76]*(15)+in_buf[77]*(17)+in_buf[78]*(6)+in_buf[79]*(17)+in_buf[80]*(-1)+in_buf[81]*(6)+in_buf[82]*(0)+in_buf[83]*(0)+in_buf[84]*(1)+in_buf[85]*(4)+in_buf[86]*(-2)+in_buf[87]*(-7)+in_buf[88]*(0)+in_buf[89]*(11)+in_buf[90]*(-10)+in_buf[91]*(7)+in_buf[92]*(41)+in_buf[93]*(26)+in_buf[94]*(32)+in_buf[95]*(7)+in_buf[96]*(13)+in_buf[97]*(1)+in_buf[98]*(11)+in_buf[99]*(5)+in_buf[100]*(-7)+in_buf[101]*(-25)+in_buf[102]*(-42)+in_buf[103]*(-39)+in_buf[104]*(-4)+in_buf[105]*(-5)+in_buf[106]*(-19)+in_buf[107]*(-15)+in_buf[108]*(15)+in_buf[109]*(16)+in_buf[110]*(6)+in_buf[111]*(-1)+in_buf[112]*(0)+in_buf[113]*(2)+in_buf[114]*(27)+in_buf[115]*(13)+in_buf[116]*(0)+in_buf[117]*(-16)+in_buf[118]*(0)+in_buf[119]*(18)+in_buf[120]*(7)+in_buf[121]*(7)+in_buf[122]*(-1)+in_buf[123]*(11)+in_buf[124]*(7)+in_buf[125]*(2)+in_buf[126]*(3)+in_buf[127]*(2)+in_buf[128]*(5)+in_buf[129]*(5)+in_buf[130]*(10)+in_buf[131]*(-4)+in_buf[132]*(11)+in_buf[133]*(22)+in_buf[134]*(14)+in_buf[135]*(-2)+in_buf[136]*(5)+in_buf[137]*(31)+in_buf[138]*(26)+in_buf[139]*(10)+in_buf[140]*(2)+in_buf[141]*(-2)+in_buf[142]*(27)+in_buf[143]*(19)+in_buf[144]*(28)+in_buf[145]*(-14)+in_buf[146]*(-11)+in_buf[147]*(12)+in_buf[148]*(13)+in_buf[149]*(5)+in_buf[150]*(2)+in_buf[151]*(1)+in_buf[152]*(-12)+in_buf[153]*(1)+in_buf[154]*(16)+in_buf[155]*(6)+in_buf[156]*(10)+in_buf[157]*(17)+in_buf[158]*(8)+in_buf[159]*(-11)+in_buf[160]*(-2)+in_buf[161]*(9)+in_buf[162]*(11)+in_buf[163]*(-1)+in_buf[164]*(-22)+in_buf[165]*(1)+in_buf[166]*(33)+in_buf[167]*(9)+in_buf[168]*(-2)+in_buf[169]*(10)+in_buf[170]*(26)+in_buf[171]*(35)+in_buf[172]*(32)+in_buf[173]*(14)+in_buf[174]*(29)+in_buf[175]*(12)+in_buf[176]*(13)+in_buf[177]*(-1)+in_buf[178]*(-10)+in_buf[179]*(0)+in_buf[180]*(-16)+in_buf[181]*(-5)+in_buf[182]*(-1)+in_buf[183]*(11)+in_buf[184]*(-1)+in_buf[185]*(0)+in_buf[186]*(1)+in_buf[187]*(-3)+in_buf[188]*(-13)+in_buf[189]*(2)+in_buf[190]*(-2)+in_buf[191]*(-5)+in_buf[192]*(6)+in_buf[193]*(3)+in_buf[194]*(12)+in_buf[195]*(27)+in_buf[196]*(-3)+in_buf[197]*(38)+in_buf[198]*(8)+in_buf[199]*(31)+in_buf[200]*(37)+in_buf[201]*(22)+in_buf[202]*(12)+in_buf[203]*(13)+in_buf[204]*(1)+in_buf[205]*(-9)+in_buf[206]*(9)+in_buf[207]*(6)+in_buf[208]*(0)+in_buf[209]*(2)+in_buf[210]*(-7)+in_buf[211]*(6)+in_buf[212]*(-1)+in_buf[213]*(4)+in_buf[214]*(18)+in_buf[215]*(4)+in_buf[216]*(0)+in_buf[217]*(0)+in_buf[218]*(0)+in_buf[219]*(-5)+in_buf[220]*(-5)+in_buf[221]*(-8)+in_buf[222]*(18)+in_buf[223]*(39)+in_buf[224]*(1)+in_buf[225]*(21)+in_buf[226]*(3)+in_buf[227]*(5)+in_buf[228]*(35)+in_buf[229]*(8)+in_buf[230]*(5)+in_buf[231]*(5)+in_buf[232]*(-1)+in_buf[233]*(0)+in_buf[234]*(12)+in_buf[235]*(14)+in_buf[236]*(18)+in_buf[237]*(22)+in_buf[238]*(17)+in_buf[239]*(3)+in_buf[240]*(13)+in_buf[241]*(15)+in_buf[242]*(22)+in_buf[243]*(5)+in_buf[244]*(14)+in_buf[245]*(5)+in_buf[246]*(17)+in_buf[247]*(17)+in_buf[248]*(7)+in_buf[249]*(-7)+in_buf[250]*(12)+in_buf[251]*(18)+in_buf[252]*(11)+in_buf[253]*(30)+in_buf[254]*(1)+in_buf[255]*(15)+in_buf[256]*(43)+in_buf[257]*(18)+in_buf[258]*(-2)+in_buf[259]*(12)+in_buf[260]*(5)+in_buf[261]*(5)+in_buf[262]*(12)+in_buf[263]*(18)+in_buf[264]*(34)+in_buf[265]*(42)+in_buf[266]*(33)+in_buf[267]*(9)+in_buf[268]*(27)+in_buf[269]*(19)+in_buf[270]*(23)+in_buf[271]*(7)+in_buf[272]*(0)+in_buf[273]*(7)+in_buf[274]*(21)+in_buf[275]*(21)+in_buf[276]*(34)+in_buf[277]*(26)+in_buf[278]*(9)+in_buf[279]*(-13)+in_buf[280]*(16)+in_buf[281]*(14)+in_buf[282]*(14)+in_buf[283]*(36)+in_buf[284]*(27)+in_buf[285]*(8)+in_buf[286]*(1)+in_buf[287]*(8)+in_buf[288]*(11)+in_buf[289]*(4)+in_buf[290]*(25)+in_buf[291]*(33)+in_buf[292]*(29)+in_buf[293]*(43)+in_buf[294]*(41)+in_buf[295]*(21)+in_buf[296]*(28)+in_buf[297]*(11)+in_buf[298]*(13)+in_buf[299]*(5)+in_buf[300]*(13)+in_buf[301]*(4)+in_buf[302]*(16)+in_buf[303]*(-13)+in_buf[304]*(25)+in_buf[305]*(36)+in_buf[306]*(44)+in_buf[307]*(-15)+in_buf[308]*(3)+in_buf[309]*(7)+in_buf[310]*(27)+in_buf[311]*(20)+in_buf[312]*(24)+in_buf[313]*(-17)+in_buf[314]*(-3)+in_buf[315]*(3)+in_buf[316]*(0)+in_buf[317]*(9)+in_buf[318]*(18)+in_buf[319]*(23)+in_buf[320]*(18)+in_buf[321]*(17)+in_buf[322]*(-10)+in_buf[323]*(-7)+in_buf[324]*(1)+in_buf[325]*(6)+in_buf[326]*(13)+in_buf[327]*(1)+in_buf[328]*(-5)+in_buf[329]*(-17)+in_buf[330]*(-12)+in_buf[331]*(-17)+in_buf[332]*(5)+in_buf[333]*(19)+in_buf[334]*(62)+in_buf[335]*(-19)+in_buf[336]*(-11)+in_buf[337]*(9)+in_buf[338]*(8)+in_buf[339]*(-9)+in_buf[340]*(-18)+in_buf[341]*(-24)+in_buf[342]*(-9)+in_buf[343]*(7)+in_buf[344]*(16)+in_buf[345]*(22)+in_buf[346]*(18)+in_buf[347]*(8)+in_buf[348]*(-3)+in_buf[349]*(-12)+in_buf[350]*(-29)+in_buf[351]*(-28)+in_buf[352]*(-17)+in_buf[353]*(-2)+in_buf[354]*(9)+in_buf[355]*(-1)+in_buf[356]*(-4)+in_buf[357]*(-15)+in_buf[358]*(-33)+in_buf[359]*(-25)+in_buf[360]*(-10)+in_buf[361]*(8)+in_buf[362]*(29)+in_buf[363]*(-36)+in_buf[364]*(2)+in_buf[365]*(9)+in_buf[366]*(0)+in_buf[367]*(-23)+in_buf[368]*(-34)+in_buf[369]*(-22)+in_buf[370]*(-7)+in_buf[371]*(-2)+in_buf[372]*(-1)+in_buf[373]*(6)+in_buf[374]*(-17)+in_buf[375]*(-19)+in_buf[376]*(-31)+in_buf[377]*(-20)+in_buf[378]*(-23)+in_buf[379]*(-21)+in_buf[380]*(-17)+in_buf[381]*(-3)+in_buf[382]*(7)+in_buf[383]*(10)+in_buf[384]*(5)+in_buf[385]*(-5)+in_buf[386]*(-16)+in_buf[387]*(-30)+in_buf[388]*(-1)+in_buf[389]*(-14)+in_buf[390]*(15)+in_buf[391]*(-2)+in_buf[392]*(16)+in_buf[393]*(7)+in_buf[394]*(10)+in_buf[395]*(-21)+in_buf[396]*(-25)+in_buf[397]*(-21)+in_buf[398]*(-29)+in_buf[399]*(-27)+in_buf[400]*(-16)+in_buf[401]*(-13)+in_buf[402]*(-30)+in_buf[403]*(-43)+in_buf[404]*(-34)+in_buf[405]*(-21)+in_buf[406]*(-10)+in_buf[407]*(-3)+in_buf[408]*(-20)+in_buf[409]*(-3)+in_buf[410]*(14)+in_buf[411]*(11)+in_buf[412]*(3)+in_buf[413]*(12)+in_buf[414]*(8)+in_buf[415]*(23)+in_buf[416]*(13)+in_buf[417]*(-26)+in_buf[418]*(-15)+in_buf[419]*(0)+in_buf[420]*(20)+in_buf[421]*(3)+in_buf[422]*(-5)+in_buf[423]*(-25)+in_buf[424]*(-16)+in_buf[425]*(-15)+in_buf[426]*(-21)+in_buf[427]*(-30)+in_buf[428]*(-20)+in_buf[429]*(-21)+in_buf[430]*(-29)+in_buf[431]*(-19)+in_buf[432]*(-5)+in_buf[433]*(-5)+in_buf[434]*(1)+in_buf[435]*(-6)+in_buf[436]*(-33)+in_buf[437]*(-17)+in_buf[438]*(4)+in_buf[439]*(7)+in_buf[440]*(26)+in_buf[441]*(30)+in_buf[442]*(35)+in_buf[443]*(37)+in_buf[444]*(34)+in_buf[445]*(-30)+in_buf[446]*(-35)+in_buf[447]*(-3)+in_buf[448]*(1)+in_buf[449]*(-2)+in_buf[450]*(3)+in_buf[451]*(0)+in_buf[452]*(0)+in_buf[453]*(-28)+in_buf[454]*(-30)+in_buf[455]*(-29)+in_buf[456]*(-19)+in_buf[457]*(-13)+in_buf[458]*(-11)+in_buf[459]*(0)+in_buf[460]*(6)+in_buf[461]*(7)+in_buf[462]*(-5)+in_buf[463]*(-16)+in_buf[464]*(-39)+in_buf[465]*(-24)+in_buf[466]*(-12)+in_buf[467]*(11)+in_buf[468]*(14)+in_buf[469]*(31)+in_buf[470]*(28)+in_buf[471]*(27)+in_buf[472]*(21)+in_buf[473]*(-41)+in_buf[474]*(-34)+in_buf[475]*(0)+in_buf[476]*(-1)+in_buf[477]*(6)+in_buf[478]*(-18)+in_buf[479]*(8)+in_buf[480]*(-10)+in_buf[481]*(-32)+in_buf[482]*(-11)+in_buf[483]*(-23)+in_buf[484]*(-14)+in_buf[485]*(-3)+in_buf[486]*(-2)+in_buf[487]*(21)+in_buf[488]*(10)+in_buf[489]*(4)+in_buf[490]*(-21)+in_buf[491]*(-28)+in_buf[492]*(-33)+in_buf[493]*(-14)+in_buf[494]*(-1)+in_buf[495]*(18)+in_buf[496]*(9)+in_buf[497]*(23)+in_buf[498]*(23)+in_buf[499]*(17)+in_buf[500]*(13)+in_buf[501]*(-10)+in_buf[502]*(-14)+in_buf[503]*(20)+in_buf[504]*(31)+in_buf[505]*(7)+in_buf[506]*(-11)+in_buf[507]*(-9)+in_buf[508]*(-24)+in_buf[509]*(-15)+in_buf[510]*(-1)+in_buf[511]*(-2)+in_buf[512]*(-2)+in_buf[513]*(-10)+in_buf[514]*(-3)+in_buf[515]*(7)+in_buf[516]*(-4)+in_buf[517]*(-33)+in_buf[518]*(-33)+in_buf[519]*(-7)+in_buf[520]*(-8)+in_buf[521]*(1)+in_buf[522]*(15)+in_buf[523]*(0)+in_buf[524]*(4)+in_buf[525]*(28)+in_buf[526]*(18)+in_buf[527]*(18)+in_buf[528]*(-8)+in_buf[529]*(-26)+in_buf[530]*(15)+in_buf[531]*(-11)+in_buf[532]*(-6)+in_buf[533]*(24)+in_buf[534]*(19)+in_buf[535]*(-1)+in_buf[536]*(-8)+in_buf[537]*(7)+in_buf[538]*(-4)+in_buf[539]*(4)+in_buf[540]*(7)+in_buf[541]*(-18)+in_buf[542]*(-15)+in_buf[543]*(-4)+in_buf[544]*(-9)+in_buf[545]*(-28)+in_buf[546]*(-24)+in_buf[547]*(-13)+in_buf[548]*(0)+in_buf[549]*(18)+in_buf[550]*(16)+in_buf[551]*(-3)+in_buf[552]*(5)+in_buf[553]*(11)+in_buf[554]*(14)+in_buf[555]*(7)+in_buf[556]*(-42)+in_buf[557]*(-46)+in_buf[558]*(13)+in_buf[559]*(-11)+in_buf[560]*(-3)+in_buf[561]*(9)+in_buf[562]*(21)+in_buf[563]*(4)+in_buf[564]*(10)+in_buf[565]*(14)+in_buf[566]*(7)+in_buf[567]*(13)+in_buf[568]*(25)+in_buf[569]*(5)+in_buf[570]*(-4)+in_buf[571]*(-6)+in_buf[572]*(-14)+in_buf[573]*(-8)+in_buf[574]*(-12)+in_buf[575]*(-1)+in_buf[576]*(17)+in_buf[577]*(24)+in_buf[578]*(11)+in_buf[579]*(10)+in_buf[580]*(-10)+in_buf[581]*(-1)+in_buf[582]*(1)+in_buf[583]*(9)+in_buf[584]*(-53)+in_buf[585]*(-38)+in_buf[586]*(3)+in_buf[587]*(-7)+in_buf[588]*(-2)+in_buf[589]*(5)+in_buf[590]*(19)+in_buf[591]*(-4)+in_buf[592]*(5)+in_buf[593]*(-2)+in_buf[594]*(-1)+in_buf[595]*(-1)+in_buf[596]*(3)+in_buf[597]*(3)+in_buf[598]*(-2)+in_buf[599]*(-2)+in_buf[600]*(-6)+in_buf[601]*(9)+in_buf[602]*(6)+in_buf[603]*(19)+in_buf[604]*(10)+in_buf[605]*(12)+in_buf[606]*(3)+in_buf[607]*(-3)+in_buf[608]*(-21)+in_buf[609]*(-16)+in_buf[610]*(13)+in_buf[611]*(-1)+in_buf[612]*(-23)+in_buf[613]*(-33)+in_buf[614]*(25)+in_buf[615]*(7)+in_buf[616]*(-1)+in_buf[617]*(8)+in_buf[618]*(14)+in_buf[619]*(22)+in_buf[620]*(-20)+in_buf[621]*(-17)+in_buf[622]*(-1)+in_buf[623]*(-6)+in_buf[624]*(-4)+in_buf[625]*(6)+in_buf[626]*(5)+in_buf[627]*(6)+in_buf[628]*(12)+in_buf[629]*(5)+in_buf[630]*(12)+in_buf[631]*(11)+in_buf[632]*(6)+in_buf[633]*(5)+in_buf[634]*(-6)+in_buf[635]*(-16)+in_buf[636]*(-17)+in_buf[637]*(-16)+in_buf[638]*(17)+in_buf[639]*(2)+in_buf[640]*(-16)+in_buf[641]*(-35)+in_buf[642]*(-17)+in_buf[643]*(7)+in_buf[644]*(-3)+in_buf[645]*(-1)+in_buf[646]*(8)+in_buf[647]*(35)+in_buf[648]*(31)+in_buf[649]*(24)+in_buf[650]*(23)+in_buf[651]*(8)+in_buf[652]*(0)+in_buf[653]*(3)+in_buf[654]*(24)+in_buf[655]*(37)+in_buf[656]*(17)+in_buf[657]*(9)+in_buf[658]*(13)+in_buf[659]*(11)+in_buf[660]*(6)+in_buf[661]*(8)+in_buf[662]*(-3)+in_buf[663]*(-3)+in_buf[664]*(-4)+in_buf[665]*(-4)+in_buf[666]*(8)+in_buf[667]*(-2)+in_buf[668]*(-7)+in_buf[669]*(-31)+in_buf[670]*(-22)+in_buf[671]*(1)+in_buf[672]*(4)+in_buf[673]*(3)+in_buf[674]*(-9)+in_buf[675]*(21)+in_buf[676]*(38)+in_buf[677]*(42)+in_buf[678]*(29)+in_buf[679]*(21)+in_buf[680]*(12)+in_buf[681]*(13)+in_buf[682]*(4)+in_buf[683]*(13)+in_buf[684]*(28)+in_buf[685]*(32)+in_buf[686]*(27)+in_buf[687]*(20)+in_buf[688]*(8)+in_buf[689]*(-1)+in_buf[690]*(11)+in_buf[691]*(8)+in_buf[692]*(-3)+in_buf[693]*(-3)+in_buf[694]*(11)+in_buf[695]*(4)+in_buf[696]*(10)+in_buf[697]*(-21)+in_buf[698]*(-23)+in_buf[699]*(0)+in_buf[700]*(0)+in_buf[701]*(2)+in_buf[702]*(-22)+in_buf[703]*(6)+in_buf[704]*(19)+in_buf[705]*(4)+in_buf[706]*(33)+in_buf[707]*(35)+in_buf[708]*(15)+in_buf[709]*(15)+in_buf[710]*(21)+in_buf[711]*(20)+in_buf[712]*(39)+in_buf[713]*(28)+in_buf[714]*(0)+in_buf[715]*(25)+in_buf[716]*(24)+in_buf[717]*(19)+in_buf[718]*(7)+in_buf[719]*(36)+in_buf[720]*(6)+in_buf[721]*(0)+in_buf[722]*(14)+in_buf[723]*(4)+in_buf[724]*(24)+in_buf[725]*(-7)+in_buf[726]*(0)+in_buf[727]*(0)+in_buf[728]*(-2)+in_buf[729]*(-1)+in_buf[730]*(0)+in_buf[731]*(19)+in_buf[732]*(-27)+in_buf[733]*(-17)+in_buf[734]*(-17)+in_buf[735]*(9)+in_buf[736]*(9)+in_buf[737]*(0)+in_buf[738]*(16)+in_buf[739]*(25)+in_buf[740]*(17)+in_buf[741]*(13)+in_buf[742]*(5)+in_buf[743]*(18)+in_buf[744]*(15)+in_buf[745]*(-2)+in_buf[746]*(-2)+in_buf[747]*(23)+in_buf[748]*(-4)+in_buf[749]*(-9)+in_buf[750]*(-13)+in_buf[751]*(9)+in_buf[752]*(-6)+in_buf[753]*(2)+in_buf[754]*(4)+in_buf[755]*(3)+in_buf[756]*(-1)+in_buf[757]*(1)+in_buf[758]*(0)+in_buf[759]*(0)+in_buf[760]*(24)+in_buf[761]*(40)+in_buf[762]*(11)+in_buf[763]*(0)+in_buf[764]*(10)+in_buf[765]*(5)+in_buf[766]*(10)+in_buf[767]*(8)+in_buf[768]*(10)+in_buf[769]*(39)+in_buf[770]*(8)+in_buf[771]*(-13)+in_buf[772]*(-1)+in_buf[773]*(23)+in_buf[774]*(3)+in_buf[775]*(-12)+in_buf[776]*(-19)+in_buf[777]*(-18)+in_buf[778]*(-12)+in_buf[779]*(23)+in_buf[780]*(2)+in_buf[781]*(-1)+in_buf[782]*(-2)+in_buf[783]*(2);
assign in_buf_weight013=in_buf[0]*(2)+in_buf[1]*(4)+in_buf[2]*(1)+in_buf[3]*(1)+in_buf[4]*(4)+in_buf[5]*(-1)+in_buf[6]*(-1)+in_buf[7]*(4)+in_buf[8]*(1)+in_buf[9]*(-3)+in_buf[10]*(1)+in_buf[11]*(-2)+in_buf[12]*(7)+in_buf[13]*(9)+in_buf[14]*(26)+in_buf[15]*(23)+in_buf[16]*(4)+in_buf[17]*(-2)+in_buf[18]*(3)+in_buf[19]*(2)+in_buf[20]*(0)+in_buf[21]*(3)+in_buf[22]*(-2)+in_buf[23]*(-3)+in_buf[24]*(0)+in_buf[25]*(3)+in_buf[26]*(0)+in_buf[27]*(0)+in_buf[28]*(-2)+in_buf[29]*(0)+in_buf[30]*(3)+in_buf[31]*(1)+in_buf[32]*(4)+in_buf[33]*(2)+in_buf[34]*(12)+in_buf[35]*(14)+in_buf[36]*(7)+in_buf[37]*(8)+in_buf[38]*(27)+in_buf[39]*(9)+in_buf[40]*(4)+in_buf[41]*(-9)+in_buf[42]*(-9)+in_buf[43]*(-6)+in_buf[44]*(-12)+in_buf[45]*(-8)+in_buf[46]*(29)+in_buf[47]*(24)+in_buf[48]*(24)+in_buf[49]*(7)+in_buf[50]*(9)+in_buf[51]*(9)+in_buf[52]*(-3)+in_buf[53]*(-1)+in_buf[54]*(0)+in_buf[55]*(2)+in_buf[56]*(0)+in_buf[57]*(2)+in_buf[58]*(18)+in_buf[59]*(7)+in_buf[60]*(15)+in_buf[61]*(9)+in_buf[62]*(7)+in_buf[63]*(10)+in_buf[64]*(34)+in_buf[65]*(57)+in_buf[66]*(59)+in_buf[67]*(60)+in_buf[68]*(45)+in_buf[69]*(28)+in_buf[70]*(44)+in_buf[71]*(69)+in_buf[72]*(49)+in_buf[73]*(34)+in_buf[74]*(31)+in_buf[75]*(24)+in_buf[76]*(35)+in_buf[77]*(48)+in_buf[78]*(32)+in_buf[79]*(28)+in_buf[80]*(22)+in_buf[81]*(3)+in_buf[82]*(-1)+in_buf[83]*(0)+in_buf[84]*(-2)+in_buf[85]*(0)+in_buf[86]*(7)+in_buf[87]*(14)+in_buf[88]*(8)+in_buf[89]*(29)+in_buf[90]*(33)+in_buf[91]*(15)+in_buf[92]*(16)+in_buf[93]*(39)+in_buf[94]*(14)+in_buf[95]*(11)+in_buf[96]*(17)+in_buf[97]*(8)+in_buf[98]*(6)+in_buf[99]*(6)+in_buf[100]*(11)+in_buf[101]*(3)+in_buf[102]*(18)+in_buf[103]*(35)+in_buf[104]*(-8)+in_buf[105]*(12)+in_buf[106]*(24)+in_buf[107]*(-2)+in_buf[108]*(3)+in_buf[109]*(-22)+in_buf[110]*(6)+in_buf[111]*(1)+in_buf[112]*(2)+in_buf[113]*(2)+in_buf[114]*(6)+in_buf[115]*(-32)+in_buf[116]*(-2)+in_buf[117]*(41)+in_buf[118]*(53)+in_buf[119]*(9)+in_buf[120]*(22)+in_buf[121]*(15)+in_buf[122]*(17)+in_buf[123]*(28)+in_buf[124]*(10)+in_buf[125]*(7)+in_buf[126]*(-8)+in_buf[127]*(-13)+in_buf[128]*(-14)+in_buf[129]*(-11)+in_buf[130]*(-2)+in_buf[131]*(23)+in_buf[132]*(8)+in_buf[133]*(-21)+in_buf[134]*(-30)+in_buf[135]*(-24)+in_buf[136]*(-12)+in_buf[137]*(-13)+in_buf[138]*(-21)+in_buf[139]*(20)+in_buf[140]*(-2)+in_buf[141]*(-1)+in_buf[142]*(42)+in_buf[143]*(0)+in_buf[144]*(19)+in_buf[145]*(36)+in_buf[146]*(39)+in_buf[147]*(11)+in_buf[148]*(13)+in_buf[149]*(-8)+in_buf[150]*(10)+in_buf[151]*(5)+in_buf[152]*(0)+in_buf[153]*(-18)+in_buf[154]*(-4)+in_buf[155]*(7)+in_buf[156]*(8)+in_buf[157]*(-7)+in_buf[158]*(-9)+in_buf[159]*(-6)+in_buf[160]*(7)+in_buf[161]*(-1)+in_buf[162]*(-19)+in_buf[163]*(4)+in_buf[164]*(5)+in_buf[165]*(-1)+in_buf[166]*(21)+in_buf[167]*(15)+in_buf[168]*(0)+in_buf[169]*(20)+in_buf[170]*(-20)+in_buf[171]*(-27)+in_buf[172]*(2)+in_buf[173]*(-13)+in_buf[174]*(-10)+in_buf[175]*(-6)+in_buf[176]*(-11)+in_buf[177]*(-14)+in_buf[178]*(-11)+in_buf[179]*(7)+in_buf[180]*(-12)+in_buf[181]*(-17)+in_buf[182]*(5)+in_buf[183]*(26)+in_buf[184]*(14)+in_buf[185]*(-14)+in_buf[186]*(-12)+in_buf[187]*(-18)+in_buf[188]*(-28)+in_buf[189]*(-24)+in_buf[190]*(-17)+in_buf[191]*(-33)+in_buf[192]*(-19)+in_buf[193]*(11)+in_buf[194]*(15)+in_buf[195]*(25)+in_buf[196]*(4)+in_buf[197]*(41)+in_buf[198]*(-12)+in_buf[199]*(-26)+in_buf[200]*(-11)+in_buf[201]*(-18)+in_buf[202]*(-21)+in_buf[203]*(0)+in_buf[204]*(-9)+in_buf[205]*(-16)+in_buf[206]*(-8)+in_buf[207]*(-2)+in_buf[208]*(-7)+in_buf[209]*(-1)+in_buf[210]*(20)+in_buf[211]*(14)+in_buf[212]*(4)+in_buf[213]*(4)+in_buf[214]*(-13)+in_buf[215]*(-25)+in_buf[216]*(-8)+in_buf[217]*(-14)+in_buf[218]*(-9)+in_buf[219]*(-45)+in_buf[220]*(-18)+in_buf[221]*(-4)+in_buf[222]*(12)+in_buf[223]*(19)+in_buf[224]*(5)+in_buf[225]*(16)+in_buf[226]*(-1)+in_buf[227]*(-32)+in_buf[228]*(-28)+in_buf[229]*(-11)+in_buf[230]*(-2)+in_buf[231]*(-4)+in_buf[232]*(-14)+in_buf[233]*(-20)+in_buf[234]*(-15)+in_buf[235]*(-20)+in_buf[236]*(-29)+in_buf[237]*(-4)+in_buf[238]*(9)+in_buf[239]*(10)+in_buf[240]*(4)+in_buf[241]*(-4)+in_buf[242]*(-30)+in_buf[243]*(-16)+in_buf[244]*(-19)+in_buf[245]*(-37)+in_buf[246]*(-37)+in_buf[247]*(-37)+in_buf[248]*(-44)+in_buf[249]*(-37)+in_buf[250]*(-17)+in_buf[251]*(-22)+in_buf[252]*(3)+in_buf[253]*(16)+in_buf[254]*(-1)+in_buf[255]*(9)+in_buf[256]*(-14)+in_buf[257]*(-3)+in_buf[258]*(-33)+in_buf[259]*(7)+in_buf[260]*(-21)+in_buf[261]*(-30)+in_buf[262]*(-31)+in_buf[263]*(-34)+in_buf[264]*(-37)+in_buf[265]*(-21)+in_buf[266]*(-4)+in_buf[267]*(29)+in_buf[268]*(13)+in_buf[269]*(-7)+in_buf[270]*(-26)+in_buf[271]*(-35)+in_buf[272]*(-37)+in_buf[273]*(-25)+in_buf[274]*(-19)+in_buf[275]*(-38)+in_buf[276]*(-29)+in_buf[277]*(-33)+in_buf[278]*(-8)+in_buf[279]*(18)+in_buf[280]*(1)+in_buf[281]*(11)+in_buf[282]*(-13)+in_buf[283]*(-37)+in_buf[284]*(-20)+in_buf[285]*(3)+in_buf[286]*(-8)+in_buf[287]*(8)+in_buf[288]*(-15)+in_buf[289]*(-22)+in_buf[290]*(-39)+in_buf[291]*(-41)+in_buf[292]*(-42)+in_buf[293]*(-22)+in_buf[294]*(9)+in_buf[295]*(34)+in_buf[296]*(18)+in_buf[297]*(0)+in_buf[298]*(-14)+in_buf[299]*(-24)+in_buf[300]*(-26)+in_buf[301]*(-4)+in_buf[302]*(0)+in_buf[303]*(-31)+in_buf[304]*(-7)+in_buf[305]*(-11)+in_buf[306]*(-9)+in_buf[307]*(5)+in_buf[308]*(0)+in_buf[309]*(9)+in_buf[310]*(-35)+in_buf[311]*(-21)+in_buf[312]*(-17)+in_buf[313]*(-2)+in_buf[314]*(-19)+in_buf[315]*(-9)+in_buf[316]*(-16)+in_buf[317]*(-29)+in_buf[318]*(-31)+in_buf[319]*(-28)+in_buf[320]*(-31)+in_buf[321]*(2)+in_buf[322]*(22)+in_buf[323]*(22)+in_buf[324]*(4)+in_buf[325]*(-14)+in_buf[326]*(-15)+in_buf[327]*(3)+in_buf[328]*(0)+in_buf[329]*(7)+in_buf[330]*(14)+in_buf[331]*(-18)+in_buf[332]*(-21)+in_buf[333]*(-12)+in_buf[334]*(-54)+in_buf[335]*(7)+in_buf[336]*(0)+in_buf[337]*(-17)+in_buf[338]*(-45)+in_buf[339]*(-4)+in_buf[340]*(-20)+in_buf[341]*(-22)+in_buf[342]*(-40)+in_buf[343]*(-7)+in_buf[344]*(-7)+in_buf[345]*(-21)+in_buf[346]*(-9)+in_buf[347]*(-10)+in_buf[348]*(11)+in_buf[349]*(20)+in_buf[350]*(36)+in_buf[351]*(8)+in_buf[352]*(-3)+in_buf[353]*(-23)+in_buf[354]*(-9)+in_buf[355]*(9)+in_buf[356]*(19)+in_buf[357]*(13)+in_buf[358]*(27)+in_buf[359]*(-2)+in_buf[360]*(5)+in_buf[361]*(7)+in_buf[362]*(-24)+in_buf[363]*(10)+in_buf[364]*(21)+in_buf[365]*(-13)+in_buf[366]*(-19)+in_buf[367]*(3)+in_buf[368]*(-17)+in_buf[369]*(-9)+in_buf[370]*(3)+in_buf[371]*(-11)+in_buf[372]*(-12)+in_buf[373]*(-2)+in_buf[374]*(13)+in_buf[375]*(21)+in_buf[376]*(35)+in_buf[377]*(26)+in_buf[378]*(24)+in_buf[379]*(10)+in_buf[380]*(3)+in_buf[381]*(-16)+in_buf[382]*(-9)+in_buf[383]*(19)+in_buf[384]*(25)+in_buf[385]*(15)+in_buf[386]*(3)+in_buf[387]*(17)+in_buf[388]*(21)+in_buf[389]*(11)+in_buf[390]*(1)+in_buf[391]*(6)+in_buf[392]*(-1)+in_buf[393]*(-15)+in_buf[394]*(-2)+in_buf[395]*(29)+in_buf[396]*(1)+in_buf[397]*(4)+in_buf[398]*(24)+in_buf[399]*(16)+in_buf[400]*(13)+in_buf[401]*(25)+in_buf[402]*(28)+in_buf[403]*(25)+in_buf[404]*(37)+in_buf[405]*(20)+in_buf[406]*(22)+in_buf[407]*(8)+in_buf[408]*(7)+in_buf[409]*(-19)+in_buf[410]*(-7)+in_buf[411]*(10)+in_buf[412]*(6)+in_buf[413]*(10)+in_buf[414]*(17)+in_buf[415]*(9)+in_buf[416]*(18)+in_buf[417]*(21)+in_buf[418]*(28)+in_buf[419]*(15)+in_buf[420]*(-2)+in_buf[421]*(-6)+in_buf[422]*(17)+in_buf[423]*(49)+in_buf[424]*(9)+in_buf[425]*(10)+in_buf[426]*(27)+in_buf[427]*(30)+in_buf[428]*(9)+in_buf[429]*(25)+in_buf[430]*(18)+in_buf[431]*(23)+in_buf[432]*(28)+in_buf[433]*(40)+in_buf[434]*(28)+in_buf[435]*(19)+in_buf[436]*(7)+in_buf[437]*(0)+in_buf[438]*(0)+in_buf[439]*(8)+in_buf[440]*(-8)+in_buf[441]*(12)+in_buf[442]*(1)+in_buf[443]*(21)+in_buf[444]*(22)+in_buf[445]*(17)+in_buf[446]*(-4)+in_buf[447]*(35)+in_buf[448]*(-2)+in_buf[449]*(-11)+in_buf[450]*(6)+in_buf[451]*(28)+in_buf[452]*(18)+in_buf[453]*(23)+in_buf[454]*(30)+in_buf[455]*(40)+in_buf[456]*(18)+in_buf[457]*(36)+in_buf[458]*(10)+in_buf[459]*(7)+in_buf[460]*(20)+in_buf[461]*(22)+in_buf[462]*(26)+in_buf[463]*(15)+in_buf[464]*(15)+in_buf[465]*(12)+in_buf[466]*(12)+in_buf[467]*(4)+in_buf[468]*(-3)+in_buf[469]*(27)+in_buf[470]*(14)+in_buf[471]*(13)+in_buf[472]*(17)+in_buf[473]*(15)+in_buf[474]*(26)+in_buf[475]*(31)+in_buf[476]*(-2)+in_buf[477]*(-1)+in_buf[478]*(22)+in_buf[479]*(23)+in_buf[480]*(12)+in_buf[481]*(24)+in_buf[482]*(31)+in_buf[483]*(13)+in_buf[484]*(12)+in_buf[485]*(16)+in_buf[486]*(18)+in_buf[487]*(8)+in_buf[488]*(8)+in_buf[489]*(15)+in_buf[490]*(20)+in_buf[491]*(10)+in_buf[492]*(14)+in_buf[493]*(8)+in_buf[494]*(9)+in_buf[495]*(0)+in_buf[496]*(9)+in_buf[497]*(19)+in_buf[498]*(29)+in_buf[499]*(15)+in_buf[500]*(6)+in_buf[501]*(22)+in_buf[502]*(18)+in_buf[503]*(-2)+in_buf[504]*(-10)+in_buf[505]*(-3)+in_buf[506]*(17)+in_buf[507]*(32)+in_buf[508]*(20)+in_buf[509]*(21)+in_buf[510]*(8)+in_buf[511]*(-3)+in_buf[512]*(5)+in_buf[513]*(8)+in_buf[514]*(-1)+in_buf[515]*(-3)+in_buf[516]*(14)+in_buf[517]*(17)+in_buf[518]*(12)+in_buf[519]*(0)+in_buf[520]*(21)+in_buf[521]*(31)+in_buf[522]*(21)+in_buf[523]*(8)+in_buf[524]*(7)+in_buf[525]*(8)+in_buf[526]*(7)+in_buf[527]*(17)+in_buf[528]*(24)+in_buf[529]*(37)+in_buf[530]*(23)+in_buf[531]*(39)+in_buf[532]*(29)+in_buf[533]*(-23)+in_buf[534]*(24)+in_buf[535]*(21)+in_buf[536]*(15)+in_buf[537]*(3)+in_buf[538]*(-3)+in_buf[539]*(0)+in_buf[540]*(-9)+in_buf[541]*(4)+in_buf[542]*(1)+in_buf[543]*(12)+in_buf[544]*(2)+in_buf[545]*(5)+in_buf[546]*(4)+in_buf[547]*(18)+in_buf[548]*(37)+in_buf[549]*(35)+in_buf[550]*(16)+in_buf[551]*(-5)+in_buf[552]*(1)+in_buf[553]*(3)+in_buf[554]*(7)+in_buf[555]*(8)+in_buf[556]*(6)+in_buf[557]*(31)+in_buf[558]*(48)+in_buf[559]*(37)+in_buf[560]*(4)+in_buf[561]*(-27)+in_buf[562]*(24)+in_buf[563]*(31)+in_buf[564]*(16)+in_buf[565]*(-3)+in_buf[566]*(2)+in_buf[567]*(6)+in_buf[568]*(-11)+in_buf[569]*(-13)+in_buf[570]*(-4)+in_buf[571]*(-2)+in_buf[572]*(-6)+in_buf[573]*(-8)+in_buf[574]*(7)+in_buf[575]*(14)+in_buf[576]*(24)+in_buf[577]*(12)+in_buf[578]*(14)+in_buf[579]*(-20)+in_buf[580]*(-9)+in_buf[581]*(-15)+in_buf[582]*(-12)+in_buf[583]*(-4)+in_buf[584]*(-15)+in_buf[585]*(-17)+in_buf[586]*(52)+in_buf[587]*(10)+in_buf[588]*(20)+in_buf[589]*(15)+in_buf[590]*(-4)+in_buf[591]*(12)+in_buf[592]*(-12)+in_buf[593]*(-19)+in_buf[594]*(-9)+in_buf[595]*(-7)+in_buf[596]*(-9)+in_buf[597]*(-4)+in_buf[598]*(-7)+in_buf[599]*(-20)+in_buf[600]*(-13)+in_buf[601]*(-18)+in_buf[602]*(1)+in_buf[603]*(-3)+in_buf[604]*(10)+in_buf[605]*(-9)+in_buf[606]*(-13)+in_buf[607]*(-25)+in_buf[608]*(-20)+in_buf[609]*(-11)+in_buf[610]*(-8)+in_buf[611]*(-26)+in_buf[612]*(-30)+in_buf[613]*(7)+in_buf[614]*(23)+in_buf[615]*(0)+in_buf[616]*(26)+in_buf[617]*(25)+in_buf[618]*(-9)+in_buf[619]*(-7)+in_buf[620]*(-42)+in_buf[621]*(-38)+in_buf[622]*(-45)+in_buf[623]*(-25)+in_buf[624]*(-19)+in_buf[625]*(-3)+in_buf[626]*(7)+in_buf[627]*(-25)+in_buf[628]*(-23)+in_buf[629]*(-25)+in_buf[630]*(-30)+in_buf[631]*(-13)+in_buf[632]*(-14)+in_buf[633]*(-28)+in_buf[634]*(-16)+in_buf[635]*(-1)+in_buf[636]*(0)+in_buf[637]*(3)+in_buf[638]*(-12)+in_buf[639]*(-52)+in_buf[640]*(-46)+in_buf[641]*(-14)+in_buf[642]*(-15)+in_buf[643]*(0)+in_buf[644]*(4)+in_buf[645]*(-1)+in_buf[646]*(11)+in_buf[647]*(-5)+in_buf[648]*(-38)+in_buf[649]*(-38)+in_buf[650]*(-22)+in_buf[651]*(-6)+in_buf[652]*(-13)+in_buf[653]*(5)+in_buf[654]*(-5)+in_buf[655]*(-3)+in_buf[656]*(4)+in_buf[657]*(-20)+in_buf[658]*(-23)+in_buf[659]*(-17)+in_buf[660]*(-21)+in_buf[661]*(-33)+in_buf[662]*(-24)+in_buf[663]*(-17)+in_buf[664]*(-9)+in_buf[665]*(11)+in_buf[666]*(-10)+in_buf[667]*(-40)+in_buf[668]*(-47)+in_buf[669]*(-9)+in_buf[670]*(10)+in_buf[671]*(5)+in_buf[672]*(-1)+in_buf[673]*(3)+in_buf[674]*(0)+in_buf[675]*(4)+in_buf[676]*(-10)+in_buf[677]*(-25)+in_buf[678]*(-25)+in_buf[679]*(-26)+in_buf[680]*(-13)+in_buf[681]*(-10)+in_buf[682]*(-6)+in_buf[683]*(7)+in_buf[684]*(0)+in_buf[685]*(-33)+in_buf[686]*(-11)+in_buf[687]*(-33)+in_buf[688]*(-14)+in_buf[689]*(-14)+in_buf[690]*(-14)+in_buf[691]*(-10)+in_buf[692]*(-1)+in_buf[693]*(33)+in_buf[694]*(-8)+in_buf[695]*(-49)+in_buf[696]*(1)+in_buf[697]*(8)+in_buf[698]*(23)+in_buf[699]*(-3)+in_buf[700]*(3)+in_buf[701]*(-1)+in_buf[702]*(3)+in_buf[703]*(3)+in_buf[704]*(2)+in_buf[705]*(-16)+in_buf[706]*(-14)+in_buf[707]*(-41)+in_buf[708]*(-60)+in_buf[709]*(-50)+in_buf[710]*(-41)+in_buf[711]*(-11)+in_buf[712]*(-15)+in_buf[713]*(-43)+in_buf[714]*(-36)+in_buf[715]*(-44)+in_buf[716]*(-44)+in_buf[717]*(-44)+in_buf[718]*(-48)+in_buf[719]*(-57)+in_buf[720]*(-15)+in_buf[721]*(-11)+in_buf[722]*(11)+in_buf[723]*(-6)+in_buf[724]*(-12)+in_buf[725]*(3)+in_buf[726]*(16)+in_buf[727]*(0)+in_buf[728]*(4)+in_buf[729]*(2)+in_buf[730]*(-1)+in_buf[731]*(-10)+in_buf[732]*(-26)+in_buf[733]*(-31)+in_buf[734]*(-34)+in_buf[735]*(-31)+in_buf[736]*(-32)+in_buf[737]*(-38)+in_buf[738]*(-46)+in_buf[739]*(-28)+in_buf[740]*(-69)+in_buf[741]*(-36)+in_buf[742]*(-70)+in_buf[743]*(-43)+in_buf[744]*(-38)+in_buf[745]*(-64)+in_buf[746]*(-74)+in_buf[747]*(-85)+in_buf[748]*(-84)+in_buf[749]*(-35)+in_buf[750]*(-30)+in_buf[751]*(-40)+in_buf[752]*(-21)+in_buf[753]*(2)+in_buf[754]*(0)+in_buf[755]*(-2)+in_buf[756]*(-2)+in_buf[757]*(3)+in_buf[758]*(-3)+in_buf[759]*(4)+in_buf[760]*(-3)+in_buf[761]*(-3)+in_buf[762]*(-15)+in_buf[763]*(-12)+in_buf[764]*(-10)+in_buf[765]*(-14)+in_buf[766]*(-28)+in_buf[767]*(-30)+in_buf[768]*(-28)+in_buf[769]*(-32)+in_buf[770]*(-44)+in_buf[771]*(-9)+in_buf[772]*(2)+in_buf[773]*(-12)+in_buf[774]*(-8)+in_buf[775]*(0)+in_buf[776]*(0)+in_buf[777]*(0)+in_buf[778]*(0)+in_buf[779]*(0)+in_buf[780]*(-1)+in_buf[781]*(-1)+in_buf[782]*(0)+in_buf[783]*(4);
assign in_buf_weight014=in_buf[0]*(0)+in_buf[1]*(1)+in_buf[2]*(-3)+in_buf[3]*(4)+in_buf[4]*(-3)+in_buf[5]*(-2)+in_buf[6]*(4)+in_buf[7]*(-3)+in_buf[8]*(0)+in_buf[9]*(3)+in_buf[10]*(2)+in_buf[11]*(2)+in_buf[12]*(3)+in_buf[13]*(3)+in_buf[14]*(7)+in_buf[15]*(6)+in_buf[16]*(0)+in_buf[17]*(4)+in_buf[18]*(4)+in_buf[19]*(3)+in_buf[20]*(3)+in_buf[21]*(-3)+in_buf[22]*(2)+in_buf[23]*(-2)+in_buf[24]*(0)+in_buf[25]*(4)+in_buf[26]*(-1)+in_buf[27]*(3)+in_buf[28]*(-3)+in_buf[29]*(4)+in_buf[30]*(-1)+in_buf[31]*(4)+in_buf[32]*(1)+in_buf[33]*(0)+in_buf[34]*(2)+in_buf[35]*(4)+in_buf[36]*(10)+in_buf[37]*(4)+in_buf[38]*(0)+in_buf[39]*(5)+in_buf[40]*(12)+in_buf[41]*(11)+in_buf[42]*(8)+in_buf[43]*(10)+in_buf[44]*(19)+in_buf[45]*(24)+in_buf[46]*(16)+in_buf[47]*(4)+in_buf[48]*(0)+in_buf[49]*(0)+in_buf[50]*(5)+in_buf[51]*(4)+in_buf[52]*(1)+in_buf[53]*(3)+in_buf[54]*(0)+in_buf[55]*(0)+in_buf[56]*(0)+in_buf[57]*(-1)+in_buf[58]*(12)+in_buf[59]*(-7)+in_buf[60]*(-2)+in_buf[61]*(1)+in_buf[62]*(7)+in_buf[63]*(5)+in_buf[64]*(9)+in_buf[65]*(35)+in_buf[66]*(48)+in_buf[67]*(21)+in_buf[68]*(22)+in_buf[69]*(6)+in_buf[70]*(8)+in_buf[71]*(26)+in_buf[72]*(20)+in_buf[73]*(15)+in_buf[74]*(6)+in_buf[75]*(-15)+in_buf[76]*(3)+in_buf[77]*(11)+in_buf[78]*(-2)+in_buf[79]*(10)+in_buf[80]*(13)+in_buf[81]*(10)+in_buf[82]*(3)+in_buf[83]*(-2)+in_buf[84]*(3)+in_buf[85]*(0)+in_buf[86]*(4)+in_buf[87]*(4)+in_buf[88]*(9)+in_buf[89]*(20)+in_buf[90]*(14)+in_buf[91]*(16)+in_buf[92]*(46)+in_buf[93]*(22)+in_buf[94]*(34)+in_buf[95]*(47)+in_buf[96]*(48)+in_buf[97]*(26)+in_buf[98]*(-3)+in_buf[99]*(29)+in_buf[100]*(28)+in_buf[101]*(23)+in_buf[102]*(48)+in_buf[103]*(38)+in_buf[104]*(13)+in_buf[105]*(22)+in_buf[106]*(15)+in_buf[107]*(23)+in_buf[108]*(28)+in_buf[109]*(-24)+in_buf[110]*(-9)+in_buf[111]*(0)+in_buf[112]*(-2)+in_buf[113]*(6)+in_buf[114]*(22)+in_buf[115]*(20)+in_buf[116]*(25)+in_buf[117]*(17)+in_buf[118]*(0)+in_buf[119]*(23)+in_buf[120]*(33)+in_buf[121]*(11)+in_buf[122]*(27)+in_buf[123]*(41)+in_buf[124]*(24)+in_buf[125]*(0)+in_buf[126]*(-3)+in_buf[127]*(1)+in_buf[128]*(8)+in_buf[129]*(16)+in_buf[130]*(33)+in_buf[131]*(35)+in_buf[132]*(18)+in_buf[133]*(-3)+in_buf[134]*(-5)+in_buf[135]*(-32)+in_buf[136]*(-15)+in_buf[137]*(-2)+in_buf[138]*(23)+in_buf[139]*(4)+in_buf[140]*(-2)+in_buf[141]*(-3)+in_buf[142]*(45)+in_buf[143]*(43)+in_buf[144]*(52)+in_buf[145]*(-5)+in_buf[146]*(-3)+in_buf[147]*(5)+in_buf[148]*(-23)+in_buf[149]*(-6)+in_buf[150]*(10)+in_buf[151]*(7)+in_buf[152]*(0)+in_buf[153]*(-10)+in_buf[154]*(-16)+in_buf[155]*(-3)+in_buf[156]*(10)+in_buf[157]*(14)+in_buf[158]*(-1)+in_buf[159]*(18)+in_buf[160]*(31)+in_buf[161]*(20)+in_buf[162]*(13)+in_buf[163]*(11)+in_buf[164]*(1)+in_buf[165]*(22)+in_buf[166]*(33)+in_buf[167]*(-7)+in_buf[168]*(-1)+in_buf[169]*(26)+in_buf[170]*(4)+in_buf[171]*(26)+in_buf[172]*(9)+in_buf[173]*(-20)+in_buf[174]*(-6)+in_buf[175]*(-9)+in_buf[176]*(-1)+in_buf[177]*(1)+in_buf[178]*(7)+in_buf[179]*(3)+in_buf[180]*(2)+in_buf[181]*(-5)+in_buf[182]*(2)+in_buf[183]*(1)+in_buf[184]*(-4)+in_buf[185]*(-10)+in_buf[186]*(-7)+in_buf[187]*(-7)+in_buf[188]*(7)+in_buf[189]*(-2)+in_buf[190]*(2)+in_buf[191]*(14)+in_buf[192]*(14)+in_buf[193]*(28)+in_buf[194]*(41)+in_buf[195]*(33)+in_buf[196]*(-11)+in_buf[197]*(23)+in_buf[198]*(-1)+in_buf[199]*(-4)+in_buf[200]*(27)+in_buf[201]*(1)+in_buf[202]*(-11)+in_buf[203]*(-8)+in_buf[204]*(20)+in_buf[205]*(3)+in_buf[206]*(-2)+in_buf[207]*(-6)+in_buf[208]*(-1)+in_buf[209]*(0)+in_buf[210]*(11)+in_buf[211]*(-5)+in_buf[212]*(-9)+in_buf[213]*(-19)+in_buf[214]*(-12)+in_buf[215]*(-2)+in_buf[216]*(-8)+in_buf[217]*(0)+in_buf[218]*(31)+in_buf[219]*(22)+in_buf[220]*(7)+in_buf[221]*(42)+in_buf[222]*(57)+in_buf[223]*(27)+in_buf[224]*(-14)+in_buf[225]*(-32)+in_buf[226]*(-6)+in_buf[227]*(15)+in_buf[228]*(19)+in_buf[229]*(-7)+in_buf[230]*(-5)+in_buf[231]*(8)+in_buf[232]*(6)+in_buf[233]*(-4)+in_buf[234]*(-8)+in_buf[235]*(-11)+in_buf[236]*(-3)+in_buf[237]*(-2)+in_buf[238]*(-1)+in_buf[239]*(-9)+in_buf[240]*(1)+in_buf[241]*(-3)+in_buf[242]*(-14)+in_buf[243]*(12)+in_buf[244]*(5)+in_buf[245]*(10)+in_buf[246]*(33)+in_buf[247]*(3)+in_buf[248]*(-4)+in_buf[249]*(41)+in_buf[250]*(55)+in_buf[251]*(12)+in_buf[252]*(-15)+in_buf[253]*(-9)+in_buf[254]*(19)+in_buf[255]*(7)+in_buf[256]*(8)+in_buf[257]*(6)+in_buf[258]*(3)+in_buf[259]*(10)+in_buf[260]*(14)+in_buf[261]*(0)+in_buf[262]*(-18)+in_buf[263]*(-20)+in_buf[264]*(-24)+in_buf[265]*(-13)+in_buf[266]*(-18)+in_buf[267]*(-9)+in_buf[268]*(10)+in_buf[269]*(-9)+in_buf[270]*(-8)+in_buf[271]*(13)+in_buf[272]*(4)+in_buf[273]*(-6)+in_buf[274]*(22)+in_buf[275]*(16)+in_buf[276]*(-17)+in_buf[277]*(27)+in_buf[278]*(53)+in_buf[279]*(12)+in_buf[280]*(-12)+in_buf[281]*(-2)+in_buf[282]*(18)+in_buf[283]*(15)+in_buf[284]*(16)+in_buf[285]*(19)+in_buf[286]*(7)+in_buf[287]*(0)+in_buf[288]*(-9)+in_buf[289]*(-29)+in_buf[290]*(-19)+in_buf[291]*(-23)+in_buf[292]*(-13)+in_buf[293]*(-8)+in_buf[294]*(-21)+in_buf[295]*(-17)+in_buf[296]*(3)+in_buf[297]*(3)+in_buf[298]*(6)+in_buf[299]*(19)+in_buf[300]*(9)+in_buf[301]*(-5)+in_buf[302]*(1)+in_buf[303]*(-4)+in_buf[304]*(-29)+in_buf[305]*(3)+in_buf[306]*(2)+in_buf[307]*(7)+in_buf[308]*(-20)+in_buf[309]*(-11)+in_buf[310]*(-31)+in_buf[311]*(17)+in_buf[312]*(35)+in_buf[313]*(-4)+in_buf[314]*(-14)+in_buf[315]*(-38)+in_buf[316]*(-38)+in_buf[317]*(-24)+in_buf[318]*(-25)+in_buf[319]*(-16)+in_buf[320]*(0)+in_buf[321]*(15)+in_buf[322]*(5)+in_buf[323]*(0)+in_buf[324]*(0)+in_buf[325]*(-5)+in_buf[326]*(-1)+in_buf[327]*(2)+in_buf[328]*(-20)+in_buf[329]*(-26)+in_buf[330]*(-41)+in_buf[331]*(-50)+in_buf[332]*(-59)+in_buf[333]*(-11)+in_buf[334]*(0)+in_buf[335]*(-10)+in_buf[336]*(-21)+in_buf[337]*(-13)+in_buf[338]*(-34)+in_buf[339]*(5)+in_buf[340]*(8)+in_buf[341]*(-19)+in_buf[342]*(-39)+in_buf[343]*(-16)+in_buf[344]*(-18)+in_buf[345]*(-5)+in_buf[346]*(3)+in_buf[347]*(9)+in_buf[348]*(25)+in_buf[349]*(16)+in_buf[350]*(13)+in_buf[351]*(3)+in_buf[352]*(0)+in_buf[353]*(0)+in_buf[354]*(-11)+in_buf[355]*(-26)+in_buf[356]*(-31)+in_buf[357]*(-44)+in_buf[358]*(-51)+in_buf[359]*(-68)+in_buf[360]*(-51)+in_buf[361]*(-21)+in_buf[362]*(1)+in_buf[363]*(-9)+in_buf[364]*(26)+in_buf[365]*(-4)+in_buf[366]*(-24)+in_buf[367]*(28)+in_buf[368]*(-16)+in_buf[369]*(-23)+in_buf[370]*(1)+in_buf[371]*(5)+in_buf[372]*(7)+in_buf[373]*(14)+in_buf[374]*(-1)+in_buf[375]*(15)+in_buf[376]*(17)+in_buf[377]*(15)+in_buf[378]*(-4)+in_buf[379]*(-1)+in_buf[380]*(0)+in_buf[381]*(-5)+in_buf[382]*(-11)+in_buf[383]*(-29)+in_buf[384]*(-37)+in_buf[385]*(-31)+in_buf[386]*(-41)+in_buf[387]*(-44)+in_buf[388]*(-43)+in_buf[389]*(-24)+in_buf[390]*(8)+in_buf[391]*(-4)+in_buf[392]*(12)+in_buf[393]*(0)+in_buf[394]*(-16)+in_buf[395]*(15)+in_buf[396]*(-24)+in_buf[397]*(-9)+in_buf[398]*(26)+in_buf[399]*(21)+in_buf[400]*(24)+in_buf[401]*(7)+in_buf[402]*(1)+in_buf[403]*(3)+in_buf[404]*(-4)+in_buf[405]*(-5)+in_buf[406]*(12)+in_buf[407]*(6)+in_buf[408]*(4)+in_buf[409]*(-11)+in_buf[410]*(-21)+in_buf[411]*(-25)+in_buf[412]*(-16)+in_buf[413]*(-2)+in_buf[414]*(-23)+in_buf[415]*(-46)+in_buf[416]*(-37)+in_buf[417]*(0)+in_buf[418]*(24)+in_buf[419]*(11)+in_buf[420]*(5)+in_buf[421]*(9)+in_buf[422]*(26)+in_buf[423]*(-1)+in_buf[424]*(-5)+in_buf[425]*(16)+in_buf[426]*(25)+in_buf[427]*(17)+in_buf[428]*(19)+in_buf[429]*(17)+in_buf[430]*(-13)+in_buf[431]*(-11)+in_buf[432]*(-9)+in_buf[433]*(4)+in_buf[434]*(17)+in_buf[435]*(-7)+in_buf[436]*(-9)+in_buf[437]*(-18)+in_buf[438]*(-23)+in_buf[439]*(-6)+in_buf[440]*(9)+in_buf[441]*(4)+in_buf[442]*(-30)+in_buf[443]*(-35)+in_buf[444]*(8)+in_buf[445]*(18)+in_buf[446]*(21)+in_buf[447]*(29)+in_buf[448]*(1)+in_buf[449]*(18)+in_buf[450]*(38)+in_buf[451]*(4)+in_buf[452]*(-7)+in_buf[453]*(4)+in_buf[454]*(2)+in_buf[455]*(3)+in_buf[456]*(-12)+in_buf[457]*(7)+in_buf[458]*(-4)+in_buf[459]*(-9)+in_buf[460]*(-12)+in_buf[461]*(14)+in_buf[462]*(2)+in_buf[463]*(-27)+in_buf[464]*(-16)+in_buf[465]*(-21)+in_buf[466]*(1)+in_buf[467]*(20)+in_buf[468]*(15)+in_buf[469]*(23)+in_buf[470]*(0)+in_buf[471]*(4)+in_buf[472]*(39)+in_buf[473]*(45)+in_buf[474]*(32)+in_buf[475]*(31)+in_buf[476]*(1)+in_buf[477]*(15)+in_buf[478]*(39)+in_buf[479]*(26)+in_buf[480]*(-9)+in_buf[481]*(-7)+in_buf[482]*(-5)+in_buf[483]*(-4)+in_buf[484]*(-7)+in_buf[485]*(-13)+in_buf[486]*(-11)+in_buf[487]*(-33)+in_buf[488]*(-16)+in_buf[489]*(2)+in_buf[490]*(-1)+in_buf[491]*(-23)+in_buf[492]*(-12)+in_buf[493]*(-11)+in_buf[494]*(-3)+in_buf[495]*(26)+in_buf[496]*(15)+in_buf[497]*(17)+in_buf[498]*(2)+in_buf[499]*(0)+in_buf[500]*(-14)+in_buf[501]*(0)+in_buf[502]*(-6)+in_buf[503]*(25)+in_buf[504]*(-33)+in_buf[505]*(18)+in_buf[506]*(34)+in_buf[507]*(19)+in_buf[508]*(-5)+in_buf[509]*(4)+in_buf[510]*(-5)+in_buf[511]*(-16)+in_buf[512]*(-16)+in_buf[513]*(-13)+in_buf[514]*(-14)+in_buf[515]*(-40)+in_buf[516]*(-22)+in_buf[517]*(4)+in_buf[518]*(4)+in_buf[519]*(-5)+in_buf[520]*(10)+in_buf[521]*(-2)+in_buf[522]*(-6)+in_buf[523]*(13)+in_buf[524]*(1)+in_buf[525]*(-6)+in_buf[526]*(-4)+in_buf[527]*(-4)+in_buf[528]*(-5)+in_buf[529]*(21)+in_buf[530]*(-13)+in_buf[531]*(35)+in_buf[532]*(26)+in_buf[533]*(-14)+in_buf[534]*(-5)+in_buf[535]*(0)+in_buf[536]*(-10)+in_buf[537]*(-3)+in_buf[538]*(-12)+in_buf[539]*(-18)+in_buf[540]*(-22)+in_buf[541]*(0)+in_buf[542]*(3)+in_buf[543]*(-17)+in_buf[544]*(-4)+in_buf[545]*(25)+in_buf[546]*(12)+in_buf[547]*(20)+in_buf[548]*(22)+in_buf[549]*(15)+in_buf[550]*(15)+in_buf[551]*(4)+in_buf[552]*(6)+in_buf[553]*(3)+in_buf[554]*(12)+in_buf[555]*(13)+in_buf[556]*(-7)+in_buf[557]*(74)+in_buf[558]*(50)+in_buf[559]*(18)+in_buf[560]*(2)+in_buf[561]*(4)+in_buf[562]*(7)+in_buf[563]*(15)+in_buf[564]*(-11)+in_buf[565]*(-14)+in_buf[566]*(-8)+in_buf[567]*(-10)+in_buf[568]*(-9)+in_buf[569]*(9)+in_buf[570]*(4)+in_buf[571]*(10)+in_buf[572]*(14)+in_buf[573]*(34)+in_buf[574]*(34)+in_buf[575]*(30)+in_buf[576]*(19)+in_buf[577]*(12)+in_buf[578]*(22)+in_buf[579]*(13)+in_buf[580]*(27)+in_buf[581]*(31)+in_buf[582]*(27)+in_buf[583]*(22)+in_buf[584]*(-11)+in_buf[585]*(50)+in_buf[586]*(35)+in_buf[587]*(5)+in_buf[588]*(0)+in_buf[589]*(15)+in_buf[590]*(19)+in_buf[591]*(34)+in_buf[592]*(-8)+in_buf[593]*(-29)+in_buf[594]*(-1)+in_buf[595]*(5)+in_buf[596]*(-1)+in_buf[597]*(8)+in_buf[598]*(7)+in_buf[599]*(25)+in_buf[600]*(24)+in_buf[601]*(30)+in_buf[602]*(26)+in_buf[603]*(13)+in_buf[604]*(10)+in_buf[605]*(13)+in_buf[606]*(27)+in_buf[607]*(34)+in_buf[608]*(11)+in_buf[609]*(13)+in_buf[610]*(33)+in_buf[611]*(34)+in_buf[612]*(5)+in_buf[613]*(34)+in_buf[614]*(31)+in_buf[615]*(1)+in_buf[616]*(-1)+in_buf[617]*(10)+in_buf[618]*(33)+in_buf[619]*(47)+in_buf[620]*(30)+in_buf[621]*(10)+in_buf[622]*(1)+in_buf[623]*(12)+in_buf[624]*(9)+in_buf[625]*(16)+in_buf[626]*(5)+in_buf[627]*(21)+in_buf[628]*(15)+in_buf[629]*(10)+in_buf[630]*(6)+in_buf[631]*(8)+in_buf[632]*(11)+in_buf[633]*(19)+in_buf[634]*(16)+in_buf[635]*(15)+in_buf[636]*(23)+in_buf[637]*(17)+in_buf[638]*(16)+in_buf[639]*(36)+in_buf[640]*(38)+in_buf[641]*(25)+in_buf[642]*(4)+in_buf[643]*(-6)+in_buf[644]*(3)+in_buf[645]*(-2)+in_buf[646]*(35)+in_buf[647]*(69)+in_buf[648]*(32)+in_buf[649]*(29)+in_buf[650]*(20)+in_buf[651]*(21)+in_buf[652]*(15)+in_buf[653]*(13)+in_buf[654]*(-1)+in_buf[655]*(9)+in_buf[656]*(3)+in_buf[657]*(-5)+in_buf[658]*(0)+in_buf[659]*(13)+in_buf[660]*(14)+in_buf[661]*(25)+in_buf[662]*(17)+in_buf[663]*(1)+in_buf[664]*(8)+in_buf[665]*(13)+in_buf[666]*(46)+in_buf[667]*(48)+in_buf[668]*(43)+in_buf[669]*(34)+in_buf[670]*(8)+in_buf[671]*(0)+in_buf[672]*(0)+in_buf[673]*(0)+in_buf[674]*(-2)+in_buf[675]*(27)+in_buf[676]*(16)+in_buf[677]*(-1)+in_buf[678]*(22)+in_buf[679]*(15)+in_buf[680]*(21)+in_buf[681]*(21)+in_buf[682]*(-13)+in_buf[683]*(-8)+in_buf[684]*(5)+in_buf[685]*(-2)+in_buf[686]*(18)+in_buf[687]*(12)+in_buf[688]*(27)+in_buf[689]*(27)+in_buf[690]*(22)+in_buf[691]*(-9)+in_buf[692]*(-22)+in_buf[693]*(-4)+in_buf[694]*(13)+in_buf[695]*(-6)+in_buf[696]*(25)+in_buf[697]*(7)+in_buf[698]*(0)+in_buf[699]*(4)+in_buf[700]*(-1)+in_buf[701]*(2)+in_buf[702]*(2)+in_buf[703]*(-12)+in_buf[704]*(-16)+in_buf[705]*(-14)+in_buf[706]*(3)+in_buf[707]*(21)+in_buf[708]*(12)+in_buf[709]*(17)+in_buf[710]*(-12)+in_buf[711]*(-32)+in_buf[712]*(14)+in_buf[713]*(6)+in_buf[714]*(0)+in_buf[715]*(2)+in_buf[716]*(12)+in_buf[717]*(20)+in_buf[718]*(19)+in_buf[719]*(12)+in_buf[720]*(-14)+in_buf[721]*(-27)+in_buf[722]*(-22)+in_buf[723]*(-23)+in_buf[724]*(6)+in_buf[725]*(0)+in_buf[726]*(6)+in_buf[727]*(4)+in_buf[728]*(1)+in_buf[729]*(0)+in_buf[730]*(2)+in_buf[731]*(-6)+in_buf[732]*(-8)+in_buf[733]*(-19)+in_buf[734]*(-40)+in_buf[735]*(-5)+in_buf[736]*(-12)+in_buf[737]*(-27)+in_buf[738]*(-27)+in_buf[739]*(-45)+in_buf[740]*(-41)+in_buf[741]*(-16)+in_buf[742]*(-33)+in_buf[743]*(-22)+in_buf[744]*(2)+in_buf[745]*(6)+in_buf[746]*(6)+in_buf[747]*(-34)+in_buf[748]*(-20)+in_buf[749]*(38)+in_buf[750]*(35)+in_buf[751]*(-3)+in_buf[752]*(-4)+in_buf[753]*(1)+in_buf[754]*(3)+in_buf[755]*(0)+in_buf[756]*(0)+in_buf[757]*(2)+in_buf[758]*(-2)+in_buf[759]*(4)+in_buf[760]*(0)+in_buf[761]*(4)+in_buf[762]*(3)+in_buf[763]*(-1)+in_buf[764]*(-3)+in_buf[765]*(1)+in_buf[766]*(-28)+in_buf[767]*(-24)+in_buf[768]*(-13)+in_buf[769]*(-20)+in_buf[770]*(-36)+in_buf[771]*(-33)+in_buf[772]*(-36)+in_buf[773]*(-44)+in_buf[774]*(-34)+in_buf[775]*(-33)+in_buf[776]*(-20)+in_buf[777]*(-3)+in_buf[778]*(-2)+in_buf[779]*(-7)+in_buf[780]*(0)+in_buf[781]*(3)+in_buf[782]*(3)+in_buf[783]*(2);
assign in_buf_weight015=in_buf[0]*(2)+in_buf[1]*(1)+in_buf[2]*(0)+in_buf[3]*(1)+in_buf[4]*(-2)+in_buf[5]*(2)+in_buf[6]*(1)+in_buf[7]*(-1)+in_buf[8]*(0)+in_buf[9]*(-2)+in_buf[10]*(4)+in_buf[11]*(-2)+in_buf[12]*(3)+in_buf[13]*(2)+in_buf[14]*(2)+in_buf[15]*(1)+in_buf[16]*(-2)+in_buf[17]*(-3)+in_buf[18]*(-2)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(2)+in_buf[22]*(-2)+in_buf[23]*(4)+in_buf[24]*(-1)+in_buf[25]*(0)+in_buf[26]*(0)+in_buf[27]*(1)+in_buf[28]*(-3)+in_buf[29]*(3)+in_buf[30]*(3)+in_buf[31]*(4)+in_buf[32]*(1)+in_buf[33]*(2)+in_buf[34]*(0)+in_buf[35]*(3)+in_buf[36]*(4)+in_buf[37]*(-3)+in_buf[38]*(1)+in_buf[39]*(-7)+in_buf[40]*(-7)+in_buf[41]*(-1)+in_buf[42]*(33)+in_buf[43]*(8)+in_buf[44]*(-34)+in_buf[45]*(-29)+in_buf[46]*(24)+in_buf[47]*(21)+in_buf[48]*(29)+in_buf[49]*(26)+in_buf[50]*(18)+in_buf[51]*(16)+in_buf[52]*(-3)+in_buf[53]*(-1)+in_buf[54]*(1)+in_buf[55]*(-1)+in_buf[56]*(3)+in_buf[57]*(2)+in_buf[58]*(1)+in_buf[59]*(2)+in_buf[60]*(10)+in_buf[61]*(0)+in_buf[62]*(1)+in_buf[63]*(-4)+in_buf[64]*(-10)+in_buf[65]*(-34)+in_buf[66]*(-40)+in_buf[67]*(-28)+in_buf[68]*(-4)+in_buf[69]*(-34)+in_buf[70]*(-2)+in_buf[71]*(7)+in_buf[72]*(15)+in_buf[73]*(62)+in_buf[74]*(35)+in_buf[75]*(58)+in_buf[76]*(51)+in_buf[77]*(26)+in_buf[78]*(31)+in_buf[79]*(30)+in_buf[80]*(6)+in_buf[81]*(-8)+in_buf[82]*(1)+in_buf[83]*(4)+in_buf[84]*(-2)+in_buf[85]*(3)+in_buf[86]*(19)+in_buf[87]*(10)+in_buf[88]*(5)+in_buf[89]*(6)+in_buf[90]*(-2)+in_buf[91]*(0)+in_buf[92]*(-23)+in_buf[93]*(-45)+in_buf[94]*(-41)+in_buf[95]*(-54)+in_buf[96]*(-62)+in_buf[97]*(-62)+in_buf[98]*(-34)+in_buf[99]*(-18)+in_buf[100]*(-22)+in_buf[101]*(0)+in_buf[102]*(8)+in_buf[103]*(-13)+in_buf[104]*(-19)+in_buf[105]*(-18)+in_buf[106]*(6)+in_buf[107]*(-2)+in_buf[108]*(-23)+in_buf[109]*(9)+in_buf[110]*(6)+in_buf[111]*(-3)+in_buf[112]*(-2)+in_buf[113]*(-1)+in_buf[114]*(19)+in_buf[115]*(11)+in_buf[116]*(-3)+in_buf[117]*(-2)+in_buf[118]*(-3)+in_buf[119]*(-32)+in_buf[120]*(-17)+in_buf[121]*(-29)+in_buf[122]*(-30)+in_buf[123]*(-37)+in_buf[124]*(-43)+in_buf[125]*(-16)+in_buf[126]*(-8)+in_buf[127]*(0)+in_buf[128]*(-9)+in_buf[129]*(-6)+in_buf[130]*(-2)+in_buf[131]*(-17)+in_buf[132]*(-17)+in_buf[133]*(-8)+in_buf[134]*(2)+in_buf[135]*(34)+in_buf[136]*(-18)+in_buf[137]*(-19)+in_buf[138]*(-9)+in_buf[139]*(2)+in_buf[140]*(4)+in_buf[141]*(2)+in_buf[142]*(17)+in_buf[143]*(-4)+in_buf[144]*(0)+in_buf[145]*(10)+in_buf[146]*(-1)+in_buf[147]*(-33)+in_buf[148]*(-47)+in_buf[149]*(-53)+in_buf[150]*(-41)+in_buf[151]*(-33)+in_buf[152]*(-20)+in_buf[153]*(-4)+in_buf[154]*(4)+in_buf[155]*(0)+in_buf[156]*(-11)+in_buf[157]*(-3)+in_buf[158]*(-7)+in_buf[159]*(-14)+in_buf[160]*(-2)+in_buf[161]*(-4)+in_buf[162]*(2)+in_buf[163]*(0)+in_buf[164]*(0)+in_buf[165]*(-13)+in_buf[166]*(0)+in_buf[167]*(22)+in_buf[168]*(0)+in_buf[169]*(-19)+in_buf[170]*(3)+in_buf[171]*(11)+in_buf[172]*(22)+in_buf[173]*(-16)+in_buf[174]*(-10)+in_buf[175]*(-12)+in_buf[176]*(-42)+in_buf[177]*(-72)+in_buf[178]*(-38)+in_buf[179]*(-21)+in_buf[180]*(-1)+in_buf[181]*(0)+in_buf[182]*(10)+in_buf[183]*(0)+in_buf[184]*(-9)+in_buf[185]*(-2)+in_buf[186]*(13)+in_buf[187]*(-4)+in_buf[188]*(-1)+in_buf[189]*(-1)+in_buf[190]*(16)+in_buf[191]*(26)+in_buf[192]*(24)+in_buf[193]*(14)+in_buf[194]*(15)+in_buf[195]*(-14)+in_buf[196]*(3)+in_buf[197]*(-34)+in_buf[198]*(3)+in_buf[199]*(6)+in_buf[200]*(7)+in_buf[201]*(-6)+in_buf[202]*(-4)+in_buf[203]*(2)+in_buf[204]*(-43)+in_buf[205]*(-47)+in_buf[206]*(-22)+in_buf[207]*(-7)+in_buf[208]*(13)+in_buf[209]*(19)+in_buf[210]*(17)+in_buf[211]*(2)+in_buf[212]*(1)+in_buf[213]*(-6)+in_buf[214]*(-6)+in_buf[215]*(-7)+in_buf[216]*(-14)+in_buf[217]*(-5)+in_buf[218]*(8)+in_buf[219]*(47)+in_buf[220]*(13)+in_buf[221]*(-5)+in_buf[222]*(14)+in_buf[223]*(-6)+in_buf[224]*(-3)+in_buf[225]*(-41)+in_buf[226]*(-4)+in_buf[227]*(-4)+in_buf[228]*(20)+in_buf[229]*(-2)+in_buf[230]*(0)+in_buf[231]*(-11)+in_buf[232]*(-36)+in_buf[233]*(-46)+in_buf[234]*(-26)+in_buf[235]*(-3)+in_buf[236]*(24)+in_buf[237]*(27)+in_buf[238]*(15)+in_buf[239]*(0)+in_buf[240]*(-8)+in_buf[241]*(-6)+in_buf[242]*(2)+in_buf[243]*(-7)+in_buf[244]*(-24)+in_buf[245]*(0)+in_buf[246]*(4)+in_buf[247]*(0)+in_buf[248]*(35)+in_buf[249]*(5)+in_buf[250]*(1)+in_buf[251]*(16)+in_buf[252]*(-2)+in_buf[253]*(-25)+in_buf[254]*(-10)+in_buf[255]*(-12)+in_buf[256]*(14)+in_buf[257]*(-18)+in_buf[258]*(-20)+in_buf[259]*(-33)+in_buf[260]*(-58)+in_buf[261]*(-52)+in_buf[262]*(-16)+in_buf[263]*(-12)+in_buf[264]*(9)+in_buf[265]*(33)+in_buf[266]*(26)+in_buf[267]*(5)+in_buf[268]*(-5)+in_buf[269]*(-11)+in_buf[270]*(0)+in_buf[271]*(4)+in_buf[272]*(-17)+in_buf[273]*(8)+in_buf[274]*(-2)+in_buf[275]*(-12)+in_buf[276]*(19)+in_buf[277]*(-2)+in_buf[278]*(15)+in_buf[279]*(-11)+in_buf[280]*(-10)+in_buf[281]*(-15)+in_buf[282]*(-18)+in_buf[283]*(-21)+in_buf[284]*(2)+in_buf[285]*(-21)+in_buf[286]*(-50)+in_buf[287]*(-46)+in_buf[288]*(-50)+in_buf[289]*(-40)+in_buf[290]*(-17)+in_buf[291]*(-10)+in_buf[292]*(18)+in_buf[293]*(27)+in_buf[294]*(31)+in_buf[295]*(25)+in_buf[296]*(-7)+in_buf[297]*(-21)+in_buf[298]*(-8)+in_buf[299]*(9)+in_buf[300]*(8)+in_buf[301]*(25)+in_buf[302]*(17)+in_buf[303]*(21)+in_buf[304]*(37)+in_buf[305]*(37)+in_buf[306]*(9)+in_buf[307]*(-21)+in_buf[308]*(-7)+in_buf[309]*(-9)+in_buf[310]*(17)+in_buf[311]*(-12)+in_buf[312]*(3)+in_buf[313]*(-4)+in_buf[314]*(-31)+in_buf[315]*(-68)+in_buf[316]*(-63)+in_buf[317]*(-40)+in_buf[318]*(-18)+in_buf[319]*(-3)+in_buf[320]*(18)+in_buf[321]*(31)+in_buf[322]*(30)+in_buf[323]*(18)+in_buf[324]*(-1)+in_buf[325]*(-6)+in_buf[326]*(-9)+in_buf[327]*(0)+in_buf[328]*(11)+in_buf[329]*(37)+in_buf[330]*(32)+in_buf[331]*(38)+in_buf[332]*(46)+in_buf[333]*(15)+in_buf[334]*(11)+in_buf[335]*(7)+in_buf[336]*(-2)+in_buf[337]*(-9)+in_buf[338]*(12)+in_buf[339]*(0)+in_buf[340]*(-1)+in_buf[341]*(-22)+in_buf[342]*(-36)+in_buf[343]*(-45)+in_buf[344]*(-47)+in_buf[345]*(-24)+in_buf[346]*(-3)+in_buf[347]*(24)+in_buf[348]*(48)+in_buf[349]*(49)+in_buf[350]*(32)+in_buf[351]*(17)+in_buf[352]*(2)+in_buf[353]*(1)+in_buf[354]*(-20)+in_buf[355]*(-10)+in_buf[356]*(23)+in_buf[357]*(42)+in_buf[358]*(10)+in_buf[359]*(21)+in_buf[360]*(22)+in_buf[361]*(-8)+in_buf[362]*(-4)+in_buf[363]*(-3)+in_buf[364]*(16)+in_buf[365]*(-3)+in_buf[366]*(-37)+in_buf[367]*(-5)+in_buf[368]*(-28)+in_buf[369]*(-51)+in_buf[370]*(-61)+in_buf[371]*(-33)+in_buf[372]*(-22)+in_buf[373]*(-5)+in_buf[374]*(-1)+in_buf[375]*(25)+in_buf[376]*(45)+in_buf[377]*(26)+in_buf[378]*(31)+in_buf[379]*(23)+in_buf[380]*(-5)+in_buf[381]*(-14)+in_buf[382]*(-37)+in_buf[383]*(-15)+in_buf[384]*(12)+in_buf[385]*(-7)+in_buf[386]*(-27)+in_buf[387]*(-22)+in_buf[388]*(-19)+in_buf[389]*(-16)+in_buf[390]*(-20)+in_buf[391]*(-4)+in_buf[392]*(7)+in_buf[393]*(1)+in_buf[394]*(-8)+in_buf[395]*(1)+in_buf[396]*(-34)+in_buf[397]*(-26)+in_buf[398]*(-54)+in_buf[399]*(-25)+in_buf[400]*(-18)+in_buf[401]*(-10)+in_buf[402]*(-6)+in_buf[403]*(12)+in_buf[404]*(26)+in_buf[405]*(32)+in_buf[406]*(34)+in_buf[407]*(15)+in_buf[408]*(-5)+in_buf[409]*(-24)+in_buf[410]*(-38)+in_buf[411]*(-20)+in_buf[412]*(-5)+in_buf[413]*(-25)+in_buf[414]*(-37)+in_buf[415]*(-33)+in_buf[416]*(-11)+in_buf[417]*(8)+in_buf[418]*(-27)+in_buf[419]*(-11)+in_buf[420]*(8)+in_buf[421]*(5)+in_buf[422]*(13)+in_buf[423]*(26)+in_buf[424]*(19)+in_buf[425]*(-17)+in_buf[426]*(-20)+in_buf[427]*(-25)+in_buf[428]*(-22)+in_buf[429]*(-15)+in_buf[430]*(-5)+in_buf[431]*(11)+in_buf[432]*(18)+in_buf[433]*(18)+in_buf[434]*(30)+in_buf[435]*(9)+in_buf[436]*(-14)+in_buf[437]*(-5)+in_buf[438]*(-8)+in_buf[439]*(-18)+in_buf[440]*(-9)+in_buf[441]*(-5)+in_buf[442]*(-16)+in_buf[443]*(-3)+in_buf[444]*(-8)+in_buf[445]*(0)+in_buf[446]*(-39)+in_buf[447]*(-18)+in_buf[448]*(-5)+in_buf[449]*(-9)+in_buf[450]*(-7)+in_buf[451]*(33)+in_buf[452]*(25)+in_buf[453]*(9)+in_buf[454]*(-24)+in_buf[455]*(-56)+in_buf[456]*(-41)+in_buf[457]*(-19)+in_buf[458]*(-16)+in_buf[459]*(2)+in_buf[460]*(16)+in_buf[461]*(26)+in_buf[462]*(27)+in_buf[463]*(2)+in_buf[464]*(-6)+in_buf[465]*(-21)+in_buf[466]*(-11)+in_buf[467]*(-18)+in_buf[468]*(-17)+in_buf[469]*(-16)+in_buf[470]*(-1)+in_buf[471]*(-1)+in_buf[472]*(-1)+in_buf[473]*(-35)+in_buf[474]*(-48)+in_buf[475]*(-13)+in_buf[476]*(-3)+in_buf[477]*(3)+in_buf[478]*(-9)+in_buf[479]*(5)+in_buf[480]*(11)+in_buf[481]*(9)+in_buf[482]*(-17)+in_buf[483]*(-30)+in_buf[484]*(-14)+in_buf[485]*(9)+in_buf[486]*(13)+in_buf[487]*(8)+in_buf[488]*(11)+in_buf[489]*(17)+in_buf[490]*(17)+in_buf[491]*(2)+in_buf[492]*(-18)+in_buf[493]*(-21)+in_buf[494]*(-4)+in_buf[495]*(-5)+in_buf[496]*(6)+in_buf[497]*(0)+in_buf[498]*(7)+in_buf[499]*(6)+in_buf[500]*(-2)+in_buf[501]*(-21)+in_buf[502]*(-34)+in_buf[503]*(-23)+in_buf[504]*(-34)+in_buf[505]*(15)+in_buf[506]*(-1)+in_buf[507]*(-22)+in_buf[508]*(-12)+in_buf[509]*(-18)+in_buf[510]*(-23)+in_buf[511]*(-6)+in_buf[512]*(-5)+in_buf[513]*(6)+in_buf[514]*(-3)+in_buf[515]*(12)+in_buf[516]*(23)+in_buf[517]*(20)+in_buf[518]*(14)+in_buf[519]*(-11)+in_buf[520]*(-25)+in_buf[521]*(-18)+in_buf[522]*(-18)+in_buf[523]*(-24)+in_buf[524]*(-10)+in_buf[525]*(-17)+in_buf[526]*(-29)+in_buf[527]*(-16)+in_buf[528]*(-1)+in_buf[529]*(8)+in_buf[530]*(24)+in_buf[531]*(8)+in_buf[532]*(20)+in_buf[533]*(-8)+in_buf[534]*(11)+in_buf[535]*(-26)+in_buf[536]*(-22)+in_buf[537]*(-25)+in_buf[538]*(-18)+in_buf[539]*(-1)+in_buf[540]*(-7)+in_buf[541]*(0)+in_buf[542]*(-12)+in_buf[543]*(0)+in_buf[544]*(13)+in_buf[545]*(3)+in_buf[546]*(-2)+in_buf[547]*(-8)+in_buf[548]*(-2)+in_buf[549]*(-15)+in_buf[550]*(-31)+in_buf[551]*(-35)+in_buf[552]*(-39)+in_buf[553]*(-32)+in_buf[554]*(-37)+in_buf[555]*(-17)+in_buf[556]*(11)+in_buf[557]*(16)+in_buf[558]*(5)+in_buf[559]*(15)+in_buf[560]*(-1)+in_buf[561]*(23)+in_buf[562]*(-7)+in_buf[563]*(-62)+in_buf[564]*(-22)+in_buf[565]*(0)+in_buf[566]*(0)+in_buf[567]*(-5)+in_buf[568]*(3)+in_buf[569]*(-9)+in_buf[570]*(0)+in_buf[571]*(0)+in_buf[572]*(5)+in_buf[573]*(-3)+in_buf[574]*(-2)+in_buf[575]*(1)+in_buf[576]*(-6)+in_buf[577]*(-5)+in_buf[578]*(-27)+in_buf[579]*(-14)+in_buf[580]*(-28)+in_buf[581]*(-39)+in_buf[582]*(-24)+in_buf[583]*(-2)+in_buf[584]*(9)+in_buf[585]*(5)+in_buf[586]*(2)+in_buf[587]*(17)+in_buf[588]*(16)+in_buf[589]*(-5)+in_buf[590]*(-18)+in_buf[591]*(-22)+in_buf[592]*(-24)+in_buf[593]*(4)+in_buf[594]*(11)+in_buf[595]*(-1)+in_buf[596]*(-3)+in_buf[597]*(-3)+in_buf[598]*(0)+in_buf[599]*(2)+in_buf[600]*(3)+in_buf[601]*(-6)+in_buf[602]*(-8)+in_buf[603]*(-8)+in_buf[604]*(-25)+in_buf[605]*(-9)+in_buf[606]*(-16)+in_buf[607]*(-26)+in_buf[608]*(-32)+in_buf[609]*(-34)+in_buf[610]*(-42)+in_buf[611]*(13)+in_buf[612]*(14)+in_buf[613]*(7)+in_buf[614]*(-20)+in_buf[615]*(1)+in_buf[616]*(14)+in_buf[617]*(6)+in_buf[618]*(-13)+in_buf[619]*(14)+in_buf[620]*(-12)+in_buf[621]*(0)+in_buf[622]*(21)+in_buf[623]*(14)+in_buf[624]*(0)+in_buf[625]*(-2)+in_buf[626]*(9)+in_buf[627]*(7)+in_buf[628]*(8)+in_buf[629]*(11)+in_buf[630]*(-2)+in_buf[631]*(-15)+in_buf[632]*(-15)+in_buf[633]*(3)+in_buf[634]*(-21)+in_buf[635]*(-25)+in_buf[636]*(-32)+in_buf[637]*(-23)+in_buf[638]*(-15)+in_buf[639]*(27)+in_buf[640]*(26)+in_buf[641]*(1)+in_buf[642]*(20)+in_buf[643]*(-1)+in_buf[644]*(-2)+in_buf[645]*(0)+in_buf[646]*(-30)+in_buf[647]*(-14)+in_buf[648]*(5)+in_buf[649]*(6)+in_buf[650]*(-2)+in_buf[651]*(8)+in_buf[652]*(27)+in_buf[653]*(29)+in_buf[654]*(11)+in_buf[655]*(3)+in_buf[656]*(22)+in_buf[657]*(22)+in_buf[658]*(13)+in_buf[659]*(-5)+in_buf[660]*(-4)+in_buf[661]*(-8)+in_buf[662]*(-31)+in_buf[663]*(-28)+in_buf[664]*(-17)+in_buf[665]*(-20)+in_buf[666]*(-10)+in_buf[667]*(6)+in_buf[668]*(-1)+in_buf[669]*(-12)+in_buf[670]*(22)+in_buf[671]*(4)+in_buf[672]*(2)+in_buf[673]*(-3)+in_buf[674]*(-11)+in_buf[675]*(-30)+in_buf[676]*(-40)+in_buf[677]*(-8)+in_buf[678]*(-23)+in_buf[679]*(1)+in_buf[680]*(9)+in_buf[681]*(13)+in_buf[682]*(8)+in_buf[683]*(6)+in_buf[684]*(7)+in_buf[685]*(6)+in_buf[686]*(-5)+in_buf[687]*(8)+in_buf[688]*(-15)+in_buf[689]*(-29)+in_buf[690]*(-24)+in_buf[691]*(-3)+in_buf[692]*(-3)+in_buf[693]*(38)+in_buf[694]*(27)+in_buf[695]*(18)+in_buf[696]*(6)+in_buf[697]*(2)+in_buf[698]*(3)+in_buf[699]*(1)+in_buf[700]*(0)+in_buf[701]*(-1)+in_buf[702]*(0)+in_buf[703]*(14)+in_buf[704]*(-21)+in_buf[705]*(-17)+in_buf[706]*(-47)+in_buf[707]*(-35)+in_buf[708]*(-30)+in_buf[709]*(-26)+in_buf[710]*(-18)+in_buf[711]*(-2)+in_buf[712]*(-5)+in_buf[713]*(-6)+in_buf[714]*(-10)+in_buf[715]*(-29)+in_buf[716]*(-44)+in_buf[717]*(-42)+in_buf[718]*(-30)+in_buf[719]*(-1)+in_buf[720]*(1)+in_buf[721]*(42)+in_buf[722]*(41)+in_buf[723]*(37)+in_buf[724]*(15)+in_buf[725]*(-3)+in_buf[726]*(-6)+in_buf[727]*(0)+in_buf[728]*(1)+in_buf[729]*(-3)+in_buf[730]*(3)+in_buf[731]*(-8)+in_buf[732]*(27)+in_buf[733]*(36)+in_buf[734]*(20)+in_buf[735]*(-3)+in_buf[736]*(1)+in_buf[737]*(11)+in_buf[738]*(-8)+in_buf[739]*(6)+in_buf[740]*(-5)+in_buf[741]*(-32)+in_buf[742]*(-13)+in_buf[743]*(-23)+in_buf[744]*(14)+in_buf[745]*(13)+in_buf[746]*(17)+in_buf[747]*(11)+in_buf[748]*(0)+in_buf[749]*(9)+in_buf[750]*(-22)+in_buf[751]*(-30)+in_buf[752]*(4)+in_buf[753]*(-8)+in_buf[754]*(-2)+in_buf[755]*(-2)+in_buf[756]*(4)+in_buf[757]*(4)+in_buf[758]*(-3)+in_buf[759]*(2)+in_buf[760]*(-19)+in_buf[761]*(-23)+in_buf[762]*(-1)+in_buf[763]*(-1)+in_buf[764]*(-4)+in_buf[765]*(13)+in_buf[766]*(26)+in_buf[767]*(19)+in_buf[768]*(2)+in_buf[769]*(0)+in_buf[770]*(34)+in_buf[771]*(15)+in_buf[772]*(6)+in_buf[773]*(18)+in_buf[774]*(22)+in_buf[775]*(1)+in_buf[776]*(-2)+in_buf[777]*(-1)+in_buf[778]*(4)+in_buf[779]*(3)+in_buf[780]*(0)+in_buf[781]*(-2)+in_buf[782]*(3)+in_buf[783]*(-2);
assign in_buf_weight016=in_buf[0]*(2)+in_buf[1]*(-3)+in_buf[2]*(4)+in_buf[3]*(2)+in_buf[4]*(3)+in_buf[5]*(2)+in_buf[6]*(-3)+in_buf[7]*(-3)+in_buf[8]*(2)+in_buf[9]*(-1)+in_buf[10]*(-3)+in_buf[11]*(2)+in_buf[12]*(1)+in_buf[13]*(-7)+in_buf[14]*(0)+in_buf[15]*(1)+in_buf[16]*(-3)+in_buf[17]*(-2)+in_buf[18]*(2)+in_buf[19]*(2)+in_buf[20]*(2)+in_buf[21]*(-2)+in_buf[22]*(-2)+in_buf[23]*(-1)+in_buf[24]*(1)+in_buf[25]*(1)+in_buf[26]*(-2)+in_buf[27]*(3)+in_buf[28]*(2)+in_buf[29]*(-2)+in_buf[30]*(2)+in_buf[31]*(-2)+in_buf[32]*(-1)+in_buf[33]*(6)+in_buf[34]*(8)+in_buf[35]*(9)+in_buf[36]*(0)+in_buf[37]*(6)+in_buf[38]*(-3)+in_buf[39]*(-11)+in_buf[40]*(-26)+in_buf[41]*(-43)+in_buf[42]*(-21)+in_buf[43]*(5)+in_buf[44]*(0)+in_buf[45]*(-2)+in_buf[46]*(0)+in_buf[47]*(12)+in_buf[48]*(5)+in_buf[49]*(-8)+in_buf[50]*(10)+in_buf[51]*(3)+in_buf[52]*(0)+in_buf[53]*(4)+in_buf[54]*(2)+in_buf[55]*(3)+in_buf[56]*(3)+in_buf[57]*(-3)+in_buf[58]*(-1)+in_buf[59]*(27)+in_buf[60]*(29)+in_buf[61]*(7)+in_buf[62]*(4)+in_buf[63]*(-3)+in_buf[64]*(3)+in_buf[65]*(4)+in_buf[66]*(19)+in_buf[67]*(-1)+in_buf[68]*(1)+in_buf[69]*(-26)+in_buf[70]*(-28)+in_buf[71]*(-30)+in_buf[72]*(-28)+in_buf[73]*(-27)+in_buf[74]*(-18)+in_buf[75]*(-12)+in_buf[76]*(-9)+in_buf[77]*(-5)+in_buf[78]*(1)+in_buf[79]*(0)+in_buf[80]*(5)+in_buf[81]*(4)+in_buf[82]*(0)+in_buf[83]*(2)+in_buf[84]*(2)+in_buf[85]*(2)+in_buf[86]*(0)+in_buf[87]*(31)+in_buf[88]*(24)+in_buf[89]*(-20)+in_buf[90]*(19)+in_buf[91]*(33)+in_buf[92]*(19)+in_buf[93]*(-13)+in_buf[94]*(-32)+in_buf[95]*(-38)+in_buf[96]*(-32)+in_buf[97]*(-31)+in_buf[98]*(-29)+in_buf[99]*(-19)+in_buf[100]*(-30)+in_buf[101]*(-52)+in_buf[102]*(0)+in_buf[103]*(0)+in_buf[104]*(-16)+in_buf[105]*(-33)+in_buf[106]*(-26)+in_buf[107]*(-13)+in_buf[108]*(-4)+in_buf[109]*(-1)+in_buf[110]*(2)+in_buf[111]*(0)+in_buf[112]*(-4)+in_buf[113]*(0)+in_buf[114]*(4)+in_buf[115]*(19)+in_buf[116]*(36)+in_buf[117]*(19)+in_buf[118]*(22)+in_buf[119]*(18)+in_buf[120]*(25)+in_buf[121]*(-13)+in_buf[122]*(-24)+in_buf[123]*(11)+in_buf[124]*(-1)+in_buf[125]*(-5)+in_buf[126]*(-10)+in_buf[127]*(-25)+in_buf[128]*(-51)+in_buf[129]*(-66)+in_buf[130]*(-56)+in_buf[131]*(-34)+in_buf[132]*(-51)+in_buf[133]*(-32)+in_buf[134]*(-36)+in_buf[135]*(-11)+in_buf[136]*(-30)+in_buf[137]*(-3)+in_buf[138]*(8)+in_buf[139]*(4)+in_buf[140]*(-1)+in_buf[141]*(0)+in_buf[142]*(5)+in_buf[143]*(29)+in_buf[144]*(21)+in_buf[145]*(24)+in_buf[146]*(13)+in_buf[147]*(15)+in_buf[148]*(16)+in_buf[149]*(-13)+in_buf[150]*(-24)+in_buf[151]*(-9)+in_buf[152]*(-16)+in_buf[153]*(-8)+in_buf[154]*(-15)+in_buf[155]*(0)+in_buf[156]*(0)+in_buf[157]*(-10)+in_buf[158]*(-2)+in_buf[159]*(-7)+in_buf[160]*(-32)+in_buf[161]*(-44)+in_buf[162]*(-31)+in_buf[163]*(-19)+in_buf[164]*(-32)+in_buf[165]*(16)+in_buf[166]*(24)+in_buf[167]*(-2)+in_buf[168]*(4)+in_buf[169]*(9)+in_buf[170]*(-9)+in_buf[171]*(30)+in_buf[172]*(26)+in_buf[173]*(-11)+in_buf[174]*(7)+in_buf[175]*(4)+in_buf[176]*(2)+in_buf[177]*(-6)+in_buf[178]*(0)+in_buf[179]*(-13)+in_buf[180]*(-13)+in_buf[181]*(-10)+in_buf[182]*(0)+in_buf[183]*(3)+in_buf[184]*(22)+in_buf[185]*(5)+in_buf[186]*(-11)+in_buf[187]*(-23)+in_buf[188]*(-7)+in_buf[189]*(0)+in_buf[190]*(-52)+in_buf[191]*(-86)+in_buf[192]*(-74)+in_buf[193]*(-32)+in_buf[194]*(-2)+in_buf[195]*(-4)+in_buf[196]*(4)+in_buf[197]*(10)+in_buf[198]*(11)+in_buf[199]*(50)+in_buf[200]*(25)+in_buf[201]*(-17)+in_buf[202]*(20)+in_buf[203]*(31)+in_buf[204]*(6)+in_buf[205]*(-8)+in_buf[206]*(-4)+in_buf[207]*(-1)+in_buf[208]*(7)+in_buf[209]*(6)+in_buf[210]*(14)+in_buf[211]*(0)+in_buf[212]*(-7)+in_buf[213]*(-12)+in_buf[214]*(-16)+in_buf[215]*(-20)+in_buf[216]*(0)+in_buf[217]*(9)+in_buf[218]*(-33)+in_buf[219]*(-53)+in_buf[220]*(-54)+in_buf[221]*(-50)+in_buf[222]*(-28)+in_buf[223]*(-19)+in_buf[224]*(-7)+in_buf[225]*(19)+in_buf[226]*(15)+in_buf[227]*(5)+in_buf[228]*(27)+in_buf[229]*(12)+in_buf[230]*(17)+in_buf[231]*(20)+in_buf[232]*(13)+in_buf[233]*(3)+in_buf[234]*(21)+in_buf[235]*(19)+in_buf[236]*(18)+in_buf[237]*(18)+in_buf[238]*(34)+in_buf[239]*(10)+in_buf[240]*(-10)+in_buf[241]*(-15)+in_buf[242]*(-13)+in_buf[243]*(-1)+in_buf[244]*(7)+in_buf[245]*(6)+in_buf[246]*(14)+in_buf[247]*(-12)+in_buf[248]*(-50)+in_buf[249]*(-65)+in_buf[250]*(-16)+in_buf[251]*(-3)+in_buf[252]*(7)+in_buf[253]*(20)+in_buf[254]*(18)+in_buf[255]*(15)+in_buf[256]*(30)+in_buf[257]*(34)+in_buf[258]*(25)+in_buf[259]*(28)+in_buf[260]*(17)+in_buf[261]*(34)+in_buf[262]*(46)+in_buf[263]*(33)+in_buf[264]*(33)+in_buf[265]*(42)+in_buf[266]*(40)+in_buf[267]*(3)+in_buf[268]*(-30)+in_buf[269]*(-10)+in_buf[270]*(-17)+in_buf[271]*(0)+in_buf[272]*(6)+in_buf[273]*(4)+in_buf[274]*(16)+in_buf[275]*(-8)+in_buf[276]*(-35)+in_buf[277]*(-29)+in_buf[278]*(13)+in_buf[279]*(27)+in_buf[280]*(12)+in_buf[281]*(14)+in_buf[282]*(8)+in_buf[283]*(3)+in_buf[284]*(-1)+in_buf[285]*(31)+in_buf[286]*(41)+in_buf[287]*(35)+in_buf[288]*(32)+in_buf[289]*(44)+in_buf[290]*(48)+in_buf[291]*(34)+in_buf[292]*(18)+in_buf[293]*(46)+in_buf[294]*(26)+in_buf[295]*(-17)+in_buf[296]*(-26)+in_buf[297]*(-15)+in_buf[298]*(-8)+in_buf[299]*(2)+in_buf[300]*(1)+in_buf[301]*(7)+in_buf[302]*(15)+in_buf[303]*(7)+in_buf[304]*(-42)+in_buf[305]*(-11)+in_buf[306]*(6)+in_buf[307]*(21)+in_buf[308]*(9)+in_buf[309]*(-3)+in_buf[310]*(31)+in_buf[311]*(15)+in_buf[312]*(32)+in_buf[313]*(45)+in_buf[314]*(27)+in_buf[315]*(27)+in_buf[316]*(20)+in_buf[317]*(30)+in_buf[318]*(16)+in_buf[319]*(9)+in_buf[320]*(-8)+in_buf[321]*(7)+in_buf[322]*(0)+in_buf[323]*(-23)+in_buf[324]*(-18)+in_buf[325]*(-1)+in_buf[326]*(8)+in_buf[327]*(-7)+in_buf[328]*(5)+in_buf[329]*(5)+in_buf[330]*(19)+in_buf[331]*(2)+in_buf[332]*(-10)+in_buf[333]*(-13)+in_buf[334]*(-48)+in_buf[335]*(24)+in_buf[336]*(17)+in_buf[337]*(17)+in_buf[338]*(17)+in_buf[339]*(6)+in_buf[340]*(30)+in_buf[341]*(19)+in_buf[342]*(-6)+in_buf[343]*(-5)+in_buf[344]*(-4)+in_buf[345]*(-15)+in_buf[346]*(-27)+in_buf[347]*(-33)+in_buf[348]*(-39)+in_buf[349]*(-35)+in_buf[350]*(-4)+in_buf[351]*(-1)+in_buf[352]*(10)+in_buf[353]*(19)+in_buf[354]*(15)+in_buf[355]*(-2)+in_buf[356]*(-7)+in_buf[357]*(-7)+in_buf[358]*(-6)+in_buf[359]*(-8)+in_buf[360]*(-34)+in_buf[361]*(2)+in_buf[362]*(-16)+in_buf[363]*(28)+in_buf[364]*(-16)+in_buf[365]*(5)+in_buf[366]*(1)+in_buf[367]*(2)+in_buf[368]*(3)+in_buf[369]*(-16)+in_buf[370]*(-30)+in_buf[371]*(-32)+in_buf[372]*(-27)+in_buf[373]*(-32)+in_buf[374]*(-39)+in_buf[375]*(-40)+in_buf[376]*(-35)+in_buf[377]*(-30)+in_buf[378]*(-2)+in_buf[379]*(-7)+in_buf[380]*(14)+in_buf[381]*(6)+in_buf[382]*(-4)+in_buf[383]*(-25)+in_buf[384]*(0)+in_buf[385]*(5)+in_buf[386]*(1)+in_buf[387]*(-4)+in_buf[388]*(8)+in_buf[389]*(17)+in_buf[390]*(7)+in_buf[391]*(6)+in_buf[392]*(-19)+in_buf[393]*(6)+in_buf[394]*(14)+in_buf[395]*(-10)+in_buf[396]*(-18)+in_buf[397]*(-45)+in_buf[398]*(-41)+in_buf[399]*(-47)+in_buf[400]*(-31)+in_buf[401]*(-30)+in_buf[402]*(-11)+in_buf[403]*(-15)+in_buf[404]*(-11)+in_buf[405]*(-7)+in_buf[406]*(-4)+in_buf[407]*(-2)+in_buf[408]*(3)+in_buf[409]*(0)+in_buf[410]*(-2)+in_buf[411]*(11)+in_buf[412]*(10)+in_buf[413]*(3)+in_buf[414]*(3)+in_buf[415]*(8)+in_buf[416]*(-21)+in_buf[417]*(-21)+in_buf[418]*(19)+in_buf[419]*(15)+in_buf[420]*(-16)+in_buf[421]*(14)+in_buf[422]*(3)+in_buf[423]*(-32)+in_buf[424]*(-46)+in_buf[425]*(-47)+in_buf[426]*(-27)+in_buf[427]*(-35)+in_buf[428]*(-11)+in_buf[429]*(-5)+in_buf[430]*(0)+in_buf[431]*(-8)+in_buf[432]*(2)+in_buf[433]*(4)+in_buf[434]*(10)+in_buf[435]*(12)+in_buf[436]*(0)+in_buf[437]*(5)+in_buf[438]*(10)+in_buf[439]*(17)+in_buf[440]*(24)+in_buf[441]*(16)+in_buf[442]*(10)+in_buf[443]*(-15)+in_buf[444]*(-5)+in_buf[445]*(-33)+in_buf[446]*(3)+in_buf[447]*(15)+in_buf[448]*(2)+in_buf[449]*(16)+in_buf[450]*(11)+in_buf[451]*(-35)+in_buf[452]*(-49)+in_buf[453]*(-45)+in_buf[454]*(-13)+in_buf[455]*(-4)+in_buf[456]*(-12)+in_buf[457]*(-12)+in_buf[458]*(-7)+in_buf[459]*(-20)+in_buf[460]*(-20)+in_buf[461]*(0)+in_buf[462]*(13)+in_buf[463]*(4)+in_buf[464]*(-2)+in_buf[465]*(8)+in_buf[466]*(10)+in_buf[467]*(23)+in_buf[468]*(17)+in_buf[469]*(26)+in_buf[470]*(-1)+in_buf[471]*(-11)+in_buf[472]*(-1)+in_buf[473]*(-33)+in_buf[474]*(34)+in_buf[475]*(14)+in_buf[476]*(0)+in_buf[477]*(13)+in_buf[478]*(7)+in_buf[479]*(-19)+in_buf[480]*(-36)+in_buf[481]*(-27)+in_buf[482]*(-21)+in_buf[483]*(-1)+in_buf[484]*(-3)+in_buf[485]*(-4)+in_buf[486]*(-14)+in_buf[487]*(-20)+in_buf[488]*(-9)+in_buf[489]*(8)+in_buf[490]*(19)+in_buf[491]*(7)+in_buf[492]*(-5)+in_buf[493]*(19)+in_buf[494]*(14)+in_buf[495]*(17)+in_buf[496]*(17)+in_buf[497]*(-4)+in_buf[498]*(-5)+in_buf[499]*(-3)+in_buf[500]*(-8)+in_buf[501]*(12)+in_buf[502]*(5)+in_buf[503]*(-12)+in_buf[504]*(4)+in_buf[505]*(4)+in_buf[506]*(18)+in_buf[507]*(3)+in_buf[508]*(-12)+in_buf[509]*(-1)+in_buf[510]*(-3)+in_buf[511]*(0)+in_buf[512]*(0)+in_buf[513]*(-8)+in_buf[514]*(-7)+in_buf[515]*(-7)+in_buf[516]*(-10)+in_buf[517]*(9)+in_buf[518]*(20)+in_buf[519]*(7)+in_buf[520]*(5)+in_buf[521]*(25)+in_buf[522]*(20)+in_buf[523]*(21)+in_buf[524]*(3)+in_buf[525]*(-13)+in_buf[526]*(10)+in_buf[527]*(-2)+in_buf[528]*(-27)+in_buf[529]*(4)+in_buf[530]*(5)+in_buf[531]*(20)+in_buf[532]*(-1)+in_buf[533]*(35)+in_buf[534]*(15)+in_buf[535]*(-12)+in_buf[536]*(17)+in_buf[537]*(15)+in_buf[538]*(-12)+in_buf[539]*(6)+in_buf[540]*(14)+in_buf[541]*(3)+in_buf[542]*(-6)+in_buf[543]*(-8)+in_buf[544]*(-10)+in_buf[545]*(1)+in_buf[546]*(20)+in_buf[547]*(14)+in_buf[548]*(11)+in_buf[549]*(7)+in_buf[550]*(1)+in_buf[551]*(14)+in_buf[552]*(-16)+in_buf[553]*(-15)+in_buf[554]*(-7)+in_buf[555]*(-21)+in_buf[556]*(-35)+in_buf[557]*(8)+in_buf[558]*(0)+in_buf[559]*(16)+in_buf[560]*(-2)+in_buf[561]*(0)+in_buf[562]*(27)+in_buf[563]*(5)+in_buf[564]*(14)+in_buf[565]*(-2)+in_buf[566]*(5)+in_buf[567]*(31)+in_buf[568]*(13)+in_buf[569]*(-11)+in_buf[570]*(-24)+in_buf[571]*(-32)+in_buf[572]*(-21)+in_buf[573]*(-4)+in_buf[574]*(22)+in_buf[575]*(7)+in_buf[576]*(5)+in_buf[577]*(-5)+in_buf[578]*(-12)+in_buf[579]*(-2)+in_buf[580]*(-21)+in_buf[581]*(-17)+in_buf[582]*(-21)+in_buf[583]*(2)+in_buf[584]*(19)+in_buf[585]*(14)+in_buf[586]*(-10)+in_buf[587]*(-3)+in_buf[588]*(1)+in_buf[589]*(24)+in_buf[590]*(30)+in_buf[591]*(7)+in_buf[592]*(13)+in_buf[593]*(0)+in_buf[594]*(-6)+in_buf[595]*(-4)+in_buf[596]*(-10)+in_buf[597]*(-25)+in_buf[598]*(-14)+in_buf[599]*(-17)+in_buf[600]*(14)+in_buf[601]*(7)+in_buf[602]*(10)+in_buf[603]*(6)+in_buf[604]*(10)+in_buf[605]*(-6)+in_buf[606]*(-8)+in_buf[607]*(-3)+in_buf[608]*(-16)+in_buf[609]*(-18)+in_buf[610]*(-13)+in_buf[611]*(2)+in_buf[612]*(19)+in_buf[613]*(9)+in_buf[614]*(-36)+in_buf[615]*(0)+in_buf[616]*(0)+in_buf[617]*(15)+in_buf[618]*(27)+in_buf[619]*(-33)+in_buf[620]*(2)+in_buf[621]*(-2)+in_buf[622]*(-10)+in_buf[623]*(-8)+in_buf[624]*(-10)+in_buf[625]*(-7)+in_buf[626]*(-13)+in_buf[627]*(-6)+in_buf[628]*(14)+in_buf[629]*(5)+in_buf[630]*(3)+in_buf[631]*(12)+in_buf[632]*(13)+in_buf[633]*(0)+in_buf[634]*(-5)+in_buf[635]*(-16)+in_buf[636]*(-14)+in_buf[637]*(-14)+in_buf[638]*(-8)+in_buf[639]*(-9)+in_buf[640]*(14)+in_buf[641]*(0)+in_buf[642]*(-40)+in_buf[643]*(-2)+in_buf[644]*(0)+in_buf[645]*(-3)+in_buf[646]*(1)+in_buf[647]*(-42)+in_buf[648]*(-16)+in_buf[649]*(-5)+in_buf[650]*(1)+in_buf[651]*(-2)+in_buf[652]*(-16)+in_buf[653]*(-12)+in_buf[654]*(-5)+in_buf[655]*(3)+in_buf[656]*(-1)+in_buf[657]*(4)+in_buf[658]*(-2)+in_buf[659]*(17)+in_buf[660]*(8)+in_buf[661]*(16)+in_buf[662]*(-8)+in_buf[663]*(-30)+in_buf[664]*(-12)+in_buf[665]*(-22)+in_buf[666]*(1)+in_buf[667]*(-5)+in_buf[668]*(0)+in_buf[669]*(-13)+in_buf[670]*(4)+in_buf[671]*(-1)+in_buf[672]*(2)+in_buf[673]*(2)+in_buf[674]*(13)+in_buf[675]*(11)+in_buf[676]*(31)+in_buf[677]*(-3)+in_buf[678]*(-30)+in_buf[679]*(-30)+in_buf[680]*(2)+in_buf[681]*(-7)+in_buf[682]*(-10)+in_buf[683]*(4)+in_buf[684]*(-21)+in_buf[685]*(-25)+in_buf[686]*(-10)+in_buf[687]*(1)+in_buf[688]*(-7)+in_buf[689]*(17)+in_buf[690]*(-10)+in_buf[691]*(-4)+in_buf[692]*(-4)+in_buf[693]*(0)+in_buf[694]*(-18)+in_buf[695]*(-1)+in_buf[696]*(17)+in_buf[697]*(6)+in_buf[698]*(21)+in_buf[699]*(4)+in_buf[700]*(2)+in_buf[701]*(-3)+in_buf[702]*(-26)+in_buf[703]*(0)+in_buf[704]*(-4)+in_buf[705]*(-11)+in_buf[706]*(-22)+in_buf[707]*(-15)+in_buf[708]*(14)+in_buf[709]*(5)+in_buf[710]*(-23)+in_buf[711]*(-19)+in_buf[712]*(3)+in_buf[713]*(-17)+in_buf[714]*(7)+in_buf[715]*(4)+in_buf[716]*(16)+in_buf[717]*(12)+in_buf[718]*(0)+in_buf[719]*(14)+in_buf[720]*(2)+in_buf[721]*(0)+in_buf[722]*(-19)+in_buf[723]*(-15)+in_buf[724]*(-4)+in_buf[725]*(4)+in_buf[726]*(16)+in_buf[727]*(2)+in_buf[728]*(0)+in_buf[729]*(-2)+in_buf[730]*(2)+in_buf[731]*(5)+in_buf[732]*(-25)+in_buf[733]*(-34)+in_buf[734]*(-30)+in_buf[735]*(2)+in_buf[736]*(11)+in_buf[737]*(30)+in_buf[738]*(30)+in_buf[739]*(16)+in_buf[740]*(3)+in_buf[741]*(22)+in_buf[742]*(39)+in_buf[743]*(19)+in_buf[744]*(16)+in_buf[745]*(25)+in_buf[746]*(41)+in_buf[747]*(63)+in_buf[748]*(52)+in_buf[749]*(27)+in_buf[750]*(5)+in_buf[751]*(-10)+in_buf[752]*(-31)+in_buf[753]*(14)+in_buf[754]*(0)+in_buf[755]*(4)+in_buf[756]*(0)+in_buf[757]*(3)+in_buf[758]*(4)+in_buf[759]*(-3)+in_buf[760]*(24)+in_buf[761]*(38)+in_buf[762]*(49)+in_buf[763]*(25)+in_buf[764]*(19)+in_buf[765]*(25)+in_buf[766]*(38)+in_buf[767]*(26)+in_buf[768]*(18)+in_buf[769]*(48)+in_buf[770]*(51)+in_buf[771]*(1)+in_buf[772]*(23)+in_buf[773]*(56)+in_buf[774]*(42)+in_buf[775]*(3)+in_buf[776]*(-5)+in_buf[777]*(25)+in_buf[778]*(14)+in_buf[779]*(24)+in_buf[780]*(-3)+in_buf[781]*(-3)+in_buf[782]*(-3)+in_buf[783]*(4);
assign in_buf_weight017=in_buf[0]*(-1)+in_buf[1]*(4)+in_buf[2]*(-1)+in_buf[3]*(0)+in_buf[4]*(-3)+in_buf[5]*(4)+in_buf[6]*(0)+in_buf[7]*(0)+in_buf[8]*(-2)+in_buf[9]*(4)+in_buf[10]*(0)+in_buf[11]*(2)+in_buf[12]*(5)+in_buf[13]*(11)+in_buf[14]*(23)+in_buf[15]*(19)+in_buf[16]*(0)+in_buf[17]*(-2)+in_buf[18]*(1)+in_buf[19]*(4)+in_buf[20]*(0)+in_buf[21]*(-2)+in_buf[22]*(4)+in_buf[23]*(0)+in_buf[24]*(-1)+in_buf[25]*(2)+in_buf[26]*(0)+in_buf[27]*(-2)+in_buf[28]*(0)+in_buf[29]*(0)+in_buf[30]*(4)+in_buf[31]*(4)+in_buf[32]*(1)+in_buf[33]*(5)+in_buf[34]*(5)+in_buf[35]*(-1)+in_buf[36]*(-2)+in_buf[37]*(-3)+in_buf[38]*(11)+in_buf[39]*(16)+in_buf[40]*(9)+in_buf[41]*(1)+in_buf[42]*(-8)+in_buf[43]*(-1)+in_buf[44]*(36)+in_buf[45]*(34)+in_buf[46]*(0)+in_buf[47]*(-20)+in_buf[48]*(-14)+in_buf[49]*(1)+in_buf[50]*(-4)+in_buf[51]*(0)+in_buf[52]*(3)+in_buf[53]*(0)+in_buf[54]*(4)+in_buf[55]*(2)+in_buf[56]*(-3)+in_buf[57]*(0)+in_buf[58]*(3)+in_buf[59]*(20)+in_buf[60]*(15)+in_buf[61]*(0)+in_buf[62]*(6)+in_buf[63]*(0)+in_buf[64]*(22)+in_buf[65]*(28)+in_buf[66]*(40)+in_buf[67]*(25)+in_buf[68]*(38)+in_buf[69]*(45)+in_buf[70]*(34)+in_buf[71]*(10)+in_buf[72]*(7)+in_buf[73]*(0)+in_buf[74]*(6)+in_buf[75]*(-22)+in_buf[76]*(-8)+in_buf[77]*(6)+in_buf[78]*(-7)+in_buf[79]*(5)+in_buf[80]*(23)+in_buf[81]*(-6)+in_buf[82]*(3)+in_buf[83]*(-2)+in_buf[84]*(-1)+in_buf[85]*(4)+in_buf[86]*(32)+in_buf[87]*(18)+in_buf[88]*(-6)+in_buf[89]*(-5)+in_buf[90]*(11)+in_buf[91]*(14)+in_buf[92]*(24)+in_buf[93]*(39)+in_buf[94]*(26)+in_buf[95]*(13)+in_buf[96]*(28)+in_buf[97]*(30)+in_buf[98]*(41)+in_buf[99]*(18)+in_buf[100]*(29)+in_buf[101]*(11)+in_buf[102]*(-5)+in_buf[103]*(-5)+in_buf[104]*(-13)+in_buf[105]*(-26)+in_buf[106]*(-29)+in_buf[107]*(-38)+in_buf[108]*(-7)+in_buf[109]*(17)+in_buf[110]*(23)+in_buf[111]*(-2)+in_buf[112]*(0)+in_buf[113]*(5)+in_buf[114]*(24)+in_buf[115]*(-26)+in_buf[116]*(-1)+in_buf[117]*(16)+in_buf[118]*(31)+in_buf[119]*(23)+in_buf[120]*(29)+in_buf[121]*(25)+in_buf[122]*(13)+in_buf[123]*(26)+in_buf[124]*(31)+in_buf[125]*(30)+in_buf[126]*(28)+in_buf[127]*(30)+in_buf[128]*(24)+in_buf[129]*(29)+in_buf[130]*(23)+in_buf[131]*(3)+in_buf[132]*(-3)+in_buf[133]*(-26)+in_buf[134]*(-18)+in_buf[135]*(-49)+in_buf[136]*(-53)+in_buf[137]*(-21)+in_buf[138]*(30)+in_buf[139]*(-3)+in_buf[140]*(1)+in_buf[141]*(-3)+in_buf[142]*(-6)+in_buf[143]*(9)+in_buf[144]*(42)+in_buf[145]*(13)+in_buf[146]*(23)+in_buf[147]*(12)+in_buf[148]*(13)+in_buf[149]*(5)+in_buf[150]*(15)+in_buf[151]*(23)+in_buf[152]*(38)+in_buf[153]*(52)+in_buf[154]*(41)+in_buf[155]*(32)+in_buf[156]*(33)+in_buf[157]*(11)+in_buf[158]*(10)+in_buf[159]*(3)+in_buf[160]*(-1)+in_buf[161]*(-14)+in_buf[162]*(1)+in_buf[163]*(-11)+in_buf[164]*(-37)+in_buf[165]*(3)+in_buf[166]*(-8)+in_buf[167]*(-7)+in_buf[168]*(2)+in_buf[169]*(18)+in_buf[170]*(27)+in_buf[171]*(7)+in_buf[172]*(17)+in_buf[173]*(3)+in_buf[174]*(16)+in_buf[175]*(-4)+in_buf[176]*(-13)+in_buf[177]*(4)+in_buf[178]*(35)+in_buf[179]*(33)+in_buf[180]*(37)+in_buf[181]*(36)+in_buf[182]*(39)+in_buf[183]*(33)+in_buf[184]*(35)+in_buf[185]*(29)+in_buf[186]*(29)+in_buf[187]*(23)+in_buf[188]*(12)+in_buf[189]*(15)+in_buf[190]*(5)+in_buf[191]*(-17)+in_buf[192]*(-39)+in_buf[193]*(-16)+in_buf[194]*(-38)+in_buf[195]*(-11)+in_buf[196]*(3)+in_buf[197]*(26)+in_buf[198]*(36)+in_buf[199]*(31)+in_buf[200]*(7)+in_buf[201]*(-24)+in_buf[202]*(-17)+in_buf[203]*(-7)+in_buf[204]*(3)+in_buf[205]*(4)+in_buf[206]*(5)+in_buf[207]*(19)+in_buf[208]*(23)+in_buf[209]*(20)+in_buf[210]*(28)+in_buf[211]*(39)+in_buf[212]*(46)+in_buf[213]*(32)+in_buf[214]*(29)+in_buf[215]*(23)+in_buf[216]*(26)+in_buf[217]*(14)+in_buf[218]*(12)+in_buf[219]*(-9)+in_buf[220]*(-21)+in_buf[221]*(-4)+in_buf[222]*(-17)+in_buf[223]*(-11)+in_buf[224]*(29)+in_buf[225]*(22)+in_buf[226]*(18)+in_buf[227]*(-16)+in_buf[228]*(-18)+in_buf[229]*(-44)+in_buf[230]*(-31)+in_buf[231]*(-14)+in_buf[232]*(10)+in_buf[233]*(-8)+in_buf[234]*(-4)+in_buf[235]*(-18)+in_buf[236]*(-25)+in_buf[237]*(-23)+in_buf[238]*(7)+in_buf[239]*(27)+in_buf[240]*(39)+in_buf[241]*(24)+in_buf[242]*(23)+in_buf[243]*(24)+in_buf[244]*(19)+in_buf[245]*(3)+in_buf[246]*(21)+in_buf[247]*(12)+in_buf[248]*(-38)+in_buf[249]*(-6)+in_buf[250]*(-29)+in_buf[251]*(-9)+in_buf[252]*(0)+in_buf[253]*(13)+in_buf[254]*(-4)+in_buf[255]*(-19)+in_buf[256]*(-27)+in_buf[257]*(-25)+in_buf[258]*(-37)+in_buf[259]*(-12)+in_buf[260]*(-8)+in_buf[261]*(-29)+in_buf[262]*(-23)+in_buf[263]*(-48)+in_buf[264]*(-40)+in_buf[265]*(-47)+in_buf[266]*(-36)+in_buf[267]*(-6)+in_buf[268]*(-1)+in_buf[269]*(13)+in_buf[270]*(16)+in_buf[271]*(25)+in_buf[272]*(6)+in_buf[273]*(-1)+in_buf[274]*(15)+in_buf[275]*(12)+in_buf[276]*(-28)+in_buf[277]*(-2)+in_buf[278]*(-24)+in_buf[279]*(10)+in_buf[280]*(0)+in_buf[281]*(-3)+in_buf[282]*(0)+in_buf[283]*(-31)+in_buf[284]*(-41)+in_buf[285]*(-32)+in_buf[286]*(-21)+in_buf[287]*(-17)+in_buf[288]*(-15)+in_buf[289]*(-45)+in_buf[290]*(-40)+in_buf[291]*(-42)+in_buf[292]*(-48)+in_buf[293]*(-49)+in_buf[294]*(-50)+in_buf[295]*(-34)+in_buf[296]*(-6)+in_buf[297]*(5)+in_buf[298]*(9)+in_buf[299]*(19)+in_buf[300]*(19)+in_buf[301]*(12)+in_buf[302]*(18)+in_buf[303]*(-13)+in_buf[304]*(-13)+in_buf[305]*(3)+in_buf[306]*(10)+in_buf[307]*(15)+in_buf[308]*(-4)+in_buf[309]*(31)+in_buf[310]*(-28)+in_buf[311]*(-49)+in_buf[312]*(-28)+in_buf[313]*(-38)+in_buf[314]*(-30)+in_buf[315]*(-14)+in_buf[316]*(-21)+in_buf[317]*(-27)+in_buf[318]*(-20)+in_buf[319]*(-14)+in_buf[320]*(-32)+in_buf[321]*(-31)+in_buf[322]*(-41)+in_buf[323]*(-39)+in_buf[324]*(-35)+in_buf[325]*(-11)+in_buf[326]*(0)+in_buf[327]*(19)+in_buf[328]*(28)+in_buf[329]*(10)+in_buf[330]*(4)+in_buf[331]*(-1)+in_buf[332]*(-13)+in_buf[333]*(-5)+in_buf[334]*(11)+in_buf[335]*(-19)+in_buf[336]*(-4)+in_buf[337]*(-20)+in_buf[338]*(-42)+in_buf[339]*(-40)+in_buf[340]*(-29)+in_buf[341]*(-32)+in_buf[342]*(-11)+in_buf[343]*(-12)+in_buf[344]*(-2)+in_buf[345]*(8)+in_buf[346]*(13)+in_buf[347]*(0)+in_buf[348]*(-7)+in_buf[349]*(-25)+in_buf[350]*(-28)+in_buf[351]*(-23)+in_buf[352]*(-24)+in_buf[353]*(-22)+in_buf[354]*(-2)+in_buf[355]*(16)+in_buf[356]*(15)+in_buf[357]*(-7)+in_buf[358]*(-15)+in_buf[359]*(0)+in_buf[360]*(-21)+in_buf[361]*(-18)+in_buf[362]*(-30)+in_buf[363]*(-27)+in_buf[364]*(-16)+in_buf[365]*(-10)+in_buf[366]*(0)+in_buf[367]*(5)+in_buf[368]*(-24)+in_buf[369]*(0)+in_buf[370]*(9)+in_buf[371]*(12)+in_buf[372]*(17)+in_buf[373]*(5)+in_buf[374]*(16)+in_buf[375]*(5)+in_buf[376]*(1)+in_buf[377]*(11)+in_buf[378]*(-5)+in_buf[379]*(-14)+in_buf[380]*(-10)+in_buf[381]*(-12)+in_buf[382]*(-7)+in_buf[383]*(9)+in_buf[384]*(1)+in_buf[385]*(-2)+in_buf[386]*(-10)+in_buf[387]*(-23)+in_buf[388]*(-15)+in_buf[389]*(-7)+in_buf[390]*(-20)+in_buf[391]*(-22)+in_buf[392]*(-23)+in_buf[393]*(-9)+in_buf[394]*(10)+in_buf[395]*(8)+in_buf[396]*(0)+in_buf[397]*(-1)+in_buf[398]*(26)+in_buf[399]*(34)+in_buf[400]*(11)+in_buf[401]*(2)+in_buf[402]*(4)+in_buf[403]*(-5)+in_buf[404]*(0)+in_buf[405]*(4)+in_buf[406]*(7)+in_buf[407]*(7)+in_buf[408]*(-9)+in_buf[409]*(-10)+in_buf[410]*(2)+in_buf[411]*(-1)+in_buf[412]*(-5)+in_buf[413]*(-7)+in_buf[414]*(5)+in_buf[415]*(-20)+in_buf[416]*(-7)+in_buf[417]*(-10)+in_buf[418]*(27)+in_buf[419]*(16)+in_buf[420]*(-17)+in_buf[421]*(-5)+in_buf[422]*(-22)+in_buf[423]*(12)+in_buf[424]*(17)+in_buf[425]*(12)+in_buf[426]*(17)+in_buf[427]*(11)+in_buf[428]*(-6)+in_buf[429]*(-6)+in_buf[430]*(-4)+in_buf[431]*(-14)+in_buf[432]*(-11)+in_buf[433]*(2)+in_buf[434]*(2)+in_buf[435]*(12)+in_buf[436]*(5)+in_buf[437]*(-9)+in_buf[438]*(-1)+in_buf[439]*(-8)+in_buf[440]*(-17)+in_buf[441]*(-3)+in_buf[442]*(-2)+in_buf[443]*(-14)+in_buf[444]*(13)+in_buf[445]*(0)+in_buf[446]*(54)+in_buf[447]*(40)+in_buf[448]*(3)+in_buf[449]*(6)+in_buf[450]*(-6)+in_buf[451]*(15)+in_buf[452]*(12)+in_buf[453]*(11)+in_buf[454]*(7)+in_buf[455]*(-9)+in_buf[456]*(-11)+in_buf[457]*(-2)+in_buf[458]*(4)+in_buf[459]*(-12)+in_buf[460]*(-6)+in_buf[461]*(5)+in_buf[462]*(-3)+in_buf[463]*(7)+in_buf[464]*(5)+in_buf[465]*(8)+in_buf[466]*(-8)+in_buf[467]*(-22)+in_buf[468]*(-23)+in_buf[469]*(-10)+in_buf[470]*(-2)+in_buf[471]*(-4)+in_buf[472]*(24)+in_buf[473]*(32)+in_buf[474]*(44)+in_buf[475]*(32)+in_buf[476]*(-1)+in_buf[477]*(-2)+in_buf[478]*(-11)+in_buf[479]*(19)+in_buf[480]*(5)+in_buf[481]*(0)+in_buf[482]*(-4)+in_buf[483]*(-16)+in_buf[484]*(-2)+in_buf[485]*(10)+in_buf[486]*(-14)+in_buf[487]*(-11)+in_buf[488]*(-15)+in_buf[489]*(-4)+in_buf[490]*(1)+in_buf[491]*(10)+in_buf[492]*(11)+in_buf[493]*(-8)+in_buf[494]*(-20)+in_buf[495]*(-12)+in_buf[496]*(-22)+in_buf[497]*(-19)+in_buf[498]*(-16)+in_buf[499]*(-29)+in_buf[500]*(-1)+in_buf[501]*(34)+in_buf[502]*(24)+in_buf[503]*(32)+in_buf[504]*(25)+in_buf[505]*(-3)+in_buf[506]*(-11)+in_buf[507]*(0)+in_buf[508]*(-2)+in_buf[509]*(-9)+in_buf[510]*(-15)+in_buf[511]*(-7)+in_buf[512]*(11)+in_buf[513]*(5)+in_buf[514]*(-1)+in_buf[515]*(-5)+in_buf[516]*(-15)+in_buf[517]*(-19)+in_buf[518]*(-10)+in_buf[519]*(4)+in_buf[520]*(18)+in_buf[521]*(10)+in_buf[522]*(0)+in_buf[523]*(-5)+in_buf[524]*(-14)+in_buf[525]*(-6)+in_buf[526]*(3)+in_buf[527]*(-6)+in_buf[528]*(7)+in_buf[529]*(41)+in_buf[530]*(36)+in_buf[531]*(34)+in_buf[532]*(-23)+in_buf[533]*(9)+in_buf[534]*(8)+in_buf[535]*(-4)+in_buf[536]*(-2)+in_buf[537]*(-3)+in_buf[538]*(-8)+in_buf[539]*(-1)+in_buf[540]*(0)+in_buf[541]*(7)+in_buf[542]*(4)+in_buf[543]*(0)+in_buf[544]*(4)+in_buf[545]*(3)+in_buf[546]*(3)+in_buf[547]*(9)+in_buf[548]*(4)+in_buf[549]*(0)+in_buf[550]*(-10)+in_buf[551]*(-9)+in_buf[552]*(-9)+in_buf[553]*(-15)+in_buf[554]*(-11)+in_buf[555]*(-23)+in_buf[556]*(-2)+in_buf[557]*(27)+in_buf[558]*(54)+in_buf[559]*(16)+in_buf[560]*(0)+in_buf[561]*(10)+in_buf[562]*(33)+in_buf[563]*(26)+in_buf[564]*(4)+in_buf[565]*(15)+in_buf[566]*(4)+in_buf[567]*(7)+in_buf[568]*(0)+in_buf[569]*(1)+in_buf[570]*(10)+in_buf[571]*(22)+in_buf[572]*(13)+in_buf[573]*(13)+in_buf[574]*(4)+in_buf[575]*(13)+in_buf[576]*(9)+in_buf[577]*(-4)+in_buf[578]*(-7)+in_buf[579]*(-4)+in_buf[580]*(-6)+in_buf[581]*(0)+in_buf[582]*(-6)+in_buf[583]*(-4)+in_buf[584]*(-15)+in_buf[585]*(-3)+in_buf[586]*(36)+in_buf[587]*(-18)+in_buf[588]*(-6)+in_buf[589]*(27)+in_buf[590]*(46)+in_buf[591]*(36)+in_buf[592]*(4)+in_buf[593]*(-1)+in_buf[594]*(-2)+in_buf[595]*(0)+in_buf[596]*(-7)+in_buf[597]*(-4)+in_buf[598]*(17)+in_buf[599]*(6)+in_buf[600]*(10)+in_buf[601]*(8)+in_buf[602]*(8)+in_buf[603]*(3)+in_buf[604]*(6)+in_buf[605]*(0)+in_buf[606]*(7)+in_buf[607]*(4)+in_buf[608]*(-1)+in_buf[609]*(16)+in_buf[610]*(23)+in_buf[611]*(20)+in_buf[612]*(1)+in_buf[613]*(3)+in_buf[614]*(30)+in_buf[615]*(3)+in_buf[616]*(-10)+in_buf[617]*(8)+in_buf[618]*(44)+in_buf[619]*(10)+in_buf[620]*(0)+in_buf[621]*(-10)+in_buf[622]*(-4)+in_buf[623]*(11)+in_buf[624]*(13)+in_buf[625]*(14)+in_buf[626]*(20)+in_buf[627]*(11)+in_buf[628]*(13)+in_buf[629]*(5)+in_buf[630]*(12)+in_buf[631]*(1)+in_buf[632]*(14)+in_buf[633]*(6)+in_buf[634]*(11)+in_buf[635]*(9)+in_buf[636]*(-5)+in_buf[637]*(-5)+in_buf[638]*(6)+in_buf[639]*(4)+in_buf[640]*(30)+in_buf[641]*(-1)+in_buf[642]*(-16)+in_buf[643]*(5)+in_buf[644]*(0)+in_buf[645]*(0)+in_buf[646]*(32)+in_buf[647]*(3)+in_buf[648]*(-12)+in_buf[649]*(-3)+in_buf[650]*(5)+in_buf[651]*(18)+in_buf[652]*(1)+in_buf[653]*(10)+in_buf[654]*(21)+in_buf[655]*(25)+in_buf[656]*(2)+in_buf[657]*(0)+in_buf[658]*(3)+in_buf[659]*(0)+in_buf[660]*(-1)+in_buf[661]*(7)+in_buf[662]*(20)+in_buf[663]*(23)+in_buf[664]*(1)+in_buf[665]*(10)+in_buf[666]*(42)+in_buf[667]*(44)+in_buf[668]*(25)+in_buf[669]*(-6)+in_buf[670]*(-23)+in_buf[671]*(4)+in_buf[672]*(2)+in_buf[673]*(-3)+in_buf[674]*(23)+in_buf[675]*(14)+in_buf[676]*(45)+in_buf[677]*(13)+in_buf[678]*(0)+in_buf[679]*(-9)+in_buf[680]*(0)+in_buf[681]*(6)+in_buf[682]*(-1)+in_buf[683]*(1)+in_buf[684]*(11)+in_buf[685]*(8)+in_buf[686]*(-1)+in_buf[687]*(3)+in_buf[688]*(-11)+in_buf[689]*(15)+in_buf[690]*(21)+in_buf[691]*(1)+in_buf[692]*(-15)+in_buf[693]*(30)+in_buf[694]*(21)+in_buf[695]*(26)+in_buf[696]*(48)+in_buf[697]*(11)+in_buf[698]*(6)+in_buf[699]*(1)+in_buf[700]*(-1)+in_buf[701]*(4)+in_buf[702]*(-26)+in_buf[703]*(13)+in_buf[704]*(30)+in_buf[705]*(5)+in_buf[706]*(7)+in_buf[707]*(6)+in_buf[708]*(17)+in_buf[709]*(30)+in_buf[710]*(15)+in_buf[711]*(25)+in_buf[712]*(19)+in_buf[713]*(-8)+in_buf[714]*(-10)+in_buf[715]*(-14)+in_buf[716]*(-20)+in_buf[717]*(-17)+in_buf[718]*(-16)+in_buf[719]*(-17)+in_buf[720]*(-4)+in_buf[721]*(9)+in_buf[722]*(-13)+in_buf[723]*(-21)+in_buf[724]*(-16)+in_buf[725]*(-10)+in_buf[726]*(5)+in_buf[727]*(-3)+in_buf[728]*(3)+in_buf[729]*(2)+in_buf[730]*(4)+in_buf[731]*(25)+in_buf[732]*(-4)+in_buf[733]*(-29)+in_buf[734]*(-24)+in_buf[735]*(19)+in_buf[736]*(36)+in_buf[737]*(38)+in_buf[738]*(35)+in_buf[739]*(23)+in_buf[740]*(0)+in_buf[741]*(0)+in_buf[742]*(17)+in_buf[743]*(10)+in_buf[744]*(26)+in_buf[745]*(15)+in_buf[746]*(-1)+in_buf[747]*(-20)+in_buf[748]*(-15)+in_buf[749]*(-8)+in_buf[750]*(9)+in_buf[751]*(19)+in_buf[752]*(-5)+in_buf[753]*(12)+in_buf[754]*(0)+in_buf[755]*(0)+in_buf[756]*(3)+in_buf[757]*(4)+in_buf[758]*(4)+in_buf[759]*(4)+in_buf[760]*(-1)+in_buf[761]*(-1)+in_buf[762]*(22)+in_buf[763]*(19)+in_buf[764]*(7)+in_buf[765]*(-14)+in_buf[766]*(17)+in_buf[767]*(23)+in_buf[768]*(19)+in_buf[769]*(7)+in_buf[770]*(-10)+in_buf[771]*(-9)+in_buf[772]*(-4)+in_buf[773]*(0)+in_buf[774]*(-2)+in_buf[775]*(-3)+in_buf[776]*(-5)+in_buf[777]*(1)+in_buf[778]*(0)+in_buf[779]*(0)+in_buf[780]*(-2)+in_buf[781]*(-2)+in_buf[782]*(0)+in_buf[783]*(0);
assign in_buf_weight018=in_buf[0]*(0)+in_buf[1]*(3)+in_buf[2]*(0)+in_buf[3]*(4)+in_buf[4]*(0)+in_buf[5]*(0)+in_buf[6]*(-1)+in_buf[7]*(2)+in_buf[8]*(1)+in_buf[9]*(0)+in_buf[10]*(0)+in_buf[11]*(-3)+in_buf[12]*(4)+in_buf[13]*(4)+in_buf[14]*(0)+in_buf[15]*(3)+in_buf[16]*(3)+in_buf[17]*(3)+in_buf[18]*(1)+in_buf[19]*(-1)+in_buf[20]*(2)+in_buf[21]*(-2)+in_buf[22]*(4)+in_buf[23]*(-3)+in_buf[24]*(0)+in_buf[25]*(2)+in_buf[26]*(4)+in_buf[27]*(1)+in_buf[28]*(0)+in_buf[29]*(-1)+in_buf[30]*(-2)+in_buf[31]*(2)+in_buf[32]*(2)+in_buf[33]*(3)+in_buf[34]*(4)+in_buf[35]*(3)+in_buf[36]*(-4)+in_buf[37]*(-6)+in_buf[38]*(-21)+in_buf[39]*(-32)+in_buf[40]*(-23)+in_buf[41]*(-19)+in_buf[42]*(26)+in_buf[43]*(13)+in_buf[44]*(-41)+in_buf[45]*(-56)+in_buf[46]*(-26)+in_buf[47]*(4)+in_buf[48]*(11)+in_buf[49]*(24)+in_buf[50]*(14)+in_buf[51]*(4)+in_buf[52]*(3)+in_buf[53]*(-3)+in_buf[54]*(2)+in_buf[55]*(4)+in_buf[56]*(3)+in_buf[57]*(-1)+in_buf[58]*(-3)+in_buf[59]*(3)+in_buf[60]*(14)+in_buf[61]*(-22)+in_buf[62]*(-17)+in_buf[63]*(-16)+in_buf[64]*(-12)+in_buf[65]*(-12)+in_buf[66]*(-41)+in_buf[67]*(-43)+in_buf[68]*(-38)+in_buf[69]*(-26)+in_buf[70]*(-21)+in_buf[71]*(4)+in_buf[72]*(14)+in_buf[73]*(7)+in_buf[74]*(9)+in_buf[75]*(22)+in_buf[76]*(10)+in_buf[77]*(-6)+in_buf[78]*(6)+in_buf[79]*(1)+in_buf[80]*(-21)+in_buf[81]*(0)+in_buf[82]*(1)+in_buf[83]*(2)+in_buf[84]*(1)+in_buf[85]*(2)+in_buf[86]*(11)+in_buf[87]*(22)+in_buf[88]*(22)+in_buf[89]*(-6)+in_buf[90]*(-2)+in_buf[91]*(-4)+in_buf[92]*(-39)+in_buf[93]*(-26)+in_buf[94]*(-12)+in_buf[95]*(-37)+in_buf[96]*(-26)+in_buf[97]*(-28)+in_buf[98]*(-13)+in_buf[99]*(9)+in_buf[100]*(14)+in_buf[101]*(37)+in_buf[102]*(25)+in_buf[103]*(6)+in_buf[104]*(24)+in_buf[105]*(-11)+in_buf[106]*(-34)+in_buf[107]*(1)+in_buf[108]*(3)+in_buf[109]*(17)+in_buf[110]*(10)+in_buf[111]*(2)+in_buf[112]*(-1)+in_buf[113]*(0)+in_buf[114]*(9)+in_buf[115]*(21)+in_buf[116]*(-4)+in_buf[117]*(-1)+in_buf[118]*(2)+in_buf[119]*(-26)+in_buf[120]*(-45)+in_buf[121]*(-45)+in_buf[122]*(-15)+in_buf[123]*(-7)+in_buf[124]*(-6)+in_buf[125]*(14)+in_buf[126]*(20)+in_buf[127]*(23)+in_buf[128]*(12)+in_buf[129]*(-4)+in_buf[130]*(-11)+in_buf[131]*(-7)+in_buf[132]*(2)+in_buf[133]*(24)+in_buf[134]*(0)+in_buf[135]*(17)+in_buf[136]*(12)+in_buf[137]*(14)+in_buf[138]*(25)+in_buf[139]*(-5)+in_buf[140]*(4)+in_buf[141]*(2)+in_buf[142]*(8)+in_buf[143]*(13)+in_buf[144]*(-22)+in_buf[145]*(1)+in_buf[146]*(-11)+in_buf[147]*(-40)+in_buf[148]*(-55)+in_buf[149]*(-45)+in_buf[150]*(-19)+in_buf[151]*(-15)+in_buf[152]*(-8)+in_buf[153]*(6)+in_buf[154]*(6)+in_buf[155]*(7)+in_buf[156]*(-5)+in_buf[157]*(3)+in_buf[158]*(-1)+in_buf[159]*(7)+in_buf[160]*(14)+in_buf[161]*(10)+in_buf[162]*(20)+in_buf[163]*(15)+in_buf[164]*(-4)+in_buf[165]*(-19)+in_buf[166]*(21)+in_buf[167]*(-1)+in_buf[168]*(0)+in_buf[169]*(-14)+in_buf[170]*(-5)+in_buf[171]*(-24)+in_buf[172]*(-27)+in_buf[173]*(-27)+in_buf[174]*(-32)+in_buf[175]*(-28)+in_buf[176]*(-23)+in_buf[177]*(-14)+in_buf[178]*(-5)+in_buf[179]*(-3)+in_buf[180]*(-2)+in_buf[181]*(8)+in_buf[182]*(2)+in_buf[183]*(2)+in_buf[184]*(-7)+in_buf[185]*(5)+in_buf[186]*(9)+in_buf[187]*(8)+in_buf[188]*(19)+in_buf[189]*(12)+in_buf[190]*(13)+in_buf[191]*(19)+in_buf[192]*(25)+in_buf[193]*(16)+in_buf[194]*(20)+in_buf[195]*(-4)+in_buf[196]*(-1)+in_buf[197]*(-12)+in_buf[198]*(-20)+in_buf[199]*(-35)+in_buf[200]*(-7)+in_buf[201]*(-8)+in_buf[202]*(-26)+in_buf[203]*(-24)+in_buf[204]*(-20)+in_buf[205]*(-18)+in_buf[206]*(-3)+in_buf[207]*(-9)+in_buf[208]*(2)+in_buf[209]*(-3)+in_buf[210]*(14)+in_buf[211]*(8)+in_buf[212]*(0)+in_buf[213]*(4)+in_buf[214]*(-12)+in_buf[215]*(-3)+in_buf[216]*(0)+in_buf[217]*(-15)+in_buf[218]*(2)+in_buf[219]*(24)+in_buf[220]*(0)+in_buf[221]*(16)+in_buf[222]*(38)+in_buf[223]*(0)+in_buf[224]*(-30)+in_buf[225]*(-41)+in_buf[226]*(-22)+in_buf[227]*(-30)+in_buf[228]*(10)+in_buf[229]*(14)+in_buf[230]*(-12)+in_buf[231]*(-20)+in_buf[232]*(-34)+in_buf[233]*(-25)+in_buf[234]*(-15)+in_buf[235]*(-12)+in_buf[236]*(2)+in_buf[237]*(5)+in_buf[238]*(8)+in_buf[239]*(1)+in_buf[240]*(-3)+in_buf[241]*(-5)+in_buf[242]*(-6)+in_buf[243]*(-15)+in_buf[244]*(-6)+in_buf[245]*(-6)+in_buf[246]*(1)+in_buf[247]*(14)+in_buf[248]*(52)+in_buf[249]*(42)+in_buf[250]*(29)+in_buf[251]*(33)+in_buf[252]*(-18)+in_buf[253]*(-20)+in_buf[254]*(-16)+in_buf[255]*(-4)+in_buf[256]*(33)+in_buf[257]*(15)+in_buf[258]*(0)+in_buf[259]*(7)+in_buf[260]*(-10)+in_buf[261]*(-12)+in_buf[262]*(-20)+in_buf[263]*(-12)+in_buf[264]*(-14)+in_buf[265]*(6)+in_buf[266]*(14)+in_buf[267]*(7)+in_buf[268]*(12)+in_buf[269]*(15)+in_buf[270]*(1)+in_buf[271]*(-3)+in_buf[272]*(4)+in_buf[273]*(2)+in_buf[274]*(11)+in_buf[275]*(38)+in_buf[276]*(57)+in_buf[277]*(53)+in_buf[278]*(25)+in_buf[279]*(-14)+in_buf[280]*(-17)+in_buf[281]*(-3)+in_buf[282]*(2)+in_buf[283]*(8)+in_buf[284]*(23)+in_buf[285]*(-14)+in_buf[286]*(-14)+in_buf[287]*(-2)+in_buf[288]*(-10)+in_buf[289]*(-37)+in_buf[290]*(-22)+in_buf[291]*(-20)+in_buf[292]*(12)+in_buf[293]*(15)+in_buf[294]*(30)+in_buf[295]*(27)+in_buf[296]*(18)+in_buf[297]*(23)+in_buf[298]*(14)+in_buf[299]*(4)+in_buf[300]*(3)+in_buf[301]*(-3)+in_buf[302]*(15)+in_buf[303]*(42)+in_buf[304]*(56)+in_buf[305]*(59)+in_buf[306]*(24)+in_buf[307]*(-15)+in_buf[308]*(-13)+in_buf[309]*(-3)+in_buf[310]*(8)+in_buf[311]*(4)+in_buf[312]*(18)+in_buf[313]*(0)+in_buf[314]*(-27)+in_buf[315]*(-11)+in_buf[316]*(-42)+in_buf[317]*(-48)+in_buf[318]*(-30)+in_buf[319]*(-18)+in_buf[320]*(0)+in_buf[321]*(9)+in_buf[322]*(15)+in_buf[323]*(12)+in_buf[324]*(22)+in_buf[325]*(27)+in_buf[326]*(32)+in_buf[327]*(7)+in_buf[328]*(-7)+in_buf[329]*(-26)+in_buf[330]*(-44)+in_buf[331]*(-19)+in_buf[332]*(5)+in_buf[333]*(19)+in_buf[334]*(2)+in_buf[335]*(22)+in_buf[336]*(-3)+in_buf[337]*(-9)+in_buf[338]*(10)+in_buf[339]*(12)+in_buf[340]*(40)+in_buf[341]*(8)+in_buf[342]*(4)+in_buf[343]*(-18)+in_buf[344]*(-46)+in_buf[345]*(-37)+in_buf[346]*(-31)+in_buf[347]*(-14)+in_buf[348]*(-4)+in_buf[349]*(5)+in_buf[350]*(16)+in_buf[351]*(13)+in_buf[352]*(10)+in_buf[353]*(21)+in_buf[354]*(22)+in_buf[355]*(20)+in_buf[356]*(-19)+in_buf[357]*(-43)+in_buf[358]*(-70)+in_buf[359]*(-80)+in_buf[360]*(-60)+in_buf[361]*(-35)+in_buf[362]*(-2)+in_buf[363]*(20)+in_buf[364]*(19)+in_buf[365]*(-13)+in_buf[366]*(-35)+in_buf[367]*(11)+in_buf[368]*(23)+in_buf[369]*(9)+in_buf[370]*(-5)+in_buf[371]*(-13)+in_buf[372]*(-30)+in_buf[373]*(-14)+in_buf[374]*(-32)+in_buf[375]*(-23)+in_buf[376]*(-10)+in_buf[377]*(-1)+in_buf[378]*(22)+in_buf[379]*(20)+in_buf[380]*(9)+in_buf[381]*(8)+in_buf[382]*(2)+in_buf[383]*(6)+in_buf[384]*(-11)+in_buf[385]*(-44)+in_buf[386]*(-87)+in_buf[387]*(-90)+in_buf[388]*(-48)+in_buf[389]*(-25)+in_buf[390]*(-4)+in_buf[391]*(1)+in_buf[392]*(4)+in_buf[393]*(-5)+in_buf[394]*(-19)+in_buf[395]*(5)+in_buf[396]*(7)+in_buf[397]*(7)+in_buf[398]*(-6)+in_buf[399]*(-16)+in_buf[400]*(-13)+in_buf[401]*(-18)+in_buf[402]*(-37)+in_buf[403]*(-22)+in_buf[404]*(1)+in_buf[405]*(23)+in_buf[406]*(31)+in_buf[407]*(24)+in_buf[408]*(8)+in_buf[409]*(-2)+in_buf[410]*(-4)+in_buf[411]*(-6)+in_buf[412]*(4)+in_buf[413]*(-23)+in_buf[414]*(-64)+in_buf[415]*(-45)+in_buf[416]*(-4)+in_buf[417]*(18)+in_buf[418]*(-7)+in_buf[419]*(0)+in_buf[420]*(6)+in_buf[421]*(6)+in_buf[422]*(3)+in_buf[423]*(-30)+in_buf[424]*(10)+in_buf[425]*(8)+in_buf[426]*(5)+in_buf[427]*(8)+in_buf[428]*(3)+in_buf[429]*(-26)+in_buf[430]*(-39)+in_buf[431]*(-32)+in_buf[432]*(0)+in_buf[433]*(13)+in_buf[434]*(12)+in_buf[435]*(-7)+in_buf[436]*(-4)+in_buf[437]*(-10)+in_buf[438]*(4)+in_buf[439]*(4)+in_buf[440]*(12)+in_buf[441]*(-7)+in_buf[442]*(-43)+in_buf[443]*(-17)+in_buf[444]*(-25)+in_buf[445]*(7)+in_buf[446]*(-14)+in_buf[447]*(-1)+in_buf[448]*(-15)+in_buf[449]*(5)+in_buf[450]*(-4)+in_buf[451]*(-8)+in_buf[452]*(45)+in_buf[453]*(22)+in_buf[454]*(3)+in_buf[455]*(11)+in_buf[456]*(-10)+in_buf[457]*(-36)+in_buf[458]*(-48)+in_buf[459]*(-37)+in_buf[460]*(-8)+in_buf[461]*(1)+in_buf[462]*(4)+in_buf[463]*(-4)+in_buf[464]*(-5)+in_buf[465]*(4)+in_buf[466]*(8)+in_buf[467]*(3)+in_buf[468]*(16)+in_buf[469]*(-16)+in_buf[470]*(-49)+in_buf[471]*(-20)+in_buf[472]*(-2)+in_buf[473]*(-16)+in_buf[474]*(-15)+in_buf[475]*(-1)+in_buf[476]*(0)+in_buf[477]*(18)+in_buf[478]*(-9)+in_buf[479]*(0)+in_buf[480]*(33)+in_buf[481]*(21)+in_buf[482]*(15)+in_buf[483]*(25)+in_buf[484]*(-3)+in_buf[485]*(-30)+in_buf[486]*(-38)+in_buf[487]*(-24)+in_buf[488]*(-19)+in_buf[489]*(-12)+in_buf[490]*(-6)+in_buf[491]*(13)+in_buf[492]*(15)+in_buf[493]*(24)+in_buf[494]*(19)+in_buf[495]*(6)+in_buf[496]*(-4)+in_buf[497]*(-33)+in_buf[498]*(-31)+in_buf[499]*(2)+in_buf[500]*(15)+in_buf[501]*(-25)+in_buf[502]*(-4)+in_buf[503]*(6)+in_buf[504]*(-29)+in_buf[505]*(12)+in_buf[506]*(-6)+in_buf[507]*(4)+in_buf[508]*(11)+in_buf[509]*(25)+in_buf[510]*(20)+in_buf[511]*(15)+in_buf[512]*(15)+in_buf[513]*(-5)+in_buf[514]*(-13)+in_buf[515]*(-4)+in_buf[516]*(-15)+in_buf[517]*(-6)+in_buf[518]*(12)+in_buf[519]*(11)+in_buf[520]*(13)+in_buf[521]*(21)+in_buf[522]*(16)+in_buf[523]*(-13)+in_buf[524]*(-26)+in_buf[525]*(-36)+in_buf[526]*(-37)+in_buf[527]*(-8)+in_buf[528]*(2)+in_buf[529]*(-17)+in_buf[530]*(7)+in_buf[531]*(10)+in_buf[532]*(17)+in_buf[533]*(-9)+in_buf[534]*(-3)+in_buf[535]*(1)+in_buf[536]*(-4)+in_buf[537]*(20)+in_buf[538]*(23)+in_buf[539]*(19)+in_buf[540]*(16)+in_buf[541]*(0)+in_buf[542]*(0)+in_buf[543]*(0)+in_buf[544]*(-2)+in_buf[545]*(-3)+in_buf[546]*(8)+in_buf[547]*(10)+in_buf[548]*(15)+in_buf[549]*(16)+in_buf[550]*(14)+in_buf[551]*(-33)+in_buf[552]*(-22)+in_buf[553]*(-25)+in_buf[554]*(-24)+in_buf[555]*(-14)+in_buf[556]*(-6)+in_buf[557]*(-3)+in_buf[558]*(4)+in_buf[559]*(7)+in_buf[560]*(-2)+in_buf[561]*(16)+in_buf[562]*(-27)+in_buf[563]*(-19)+in_buf[564]*(6)+in_buf[565]*(13)+in_buf[566]*(23)+in_buf[567]*(2)+in_buf[568]*(9)+in_buf[569]*(-4)+in_buf[570]*(2)+in_buf[571]*(10)+in_buf[572]*(4)+in_buf[573]*(2)+in_buf[574]*(12)+in_buf[575]*(14)+in_buf[576]*(15)+in_buf[577]*(22)+in_buf[578]*(-1)+in_buf[579]*(-26)+in_buf[580]*(-28)+in_buf[581]*(-19)+in_buf[582]*(-16)+in_buf[583]*(-33)+in_buf[584]*(-55)+in_buf[585]*(-41)+in_buf[586]*(1)+in_buf[587]*(13)+in_buf[588]*(-3)+in_buf[589]*(-8)+in_buf[590]*(-30)+in_buf[591]*(-22)+in_buf[592]*(-13)+in_buf[593]*(4)+in_buf[594]*(22)+in_buf[595]*(17)+in_buf[596]*(2)+in_buf[597]*(-9)+in_buf[598]*(-1)+in_buf[599]*(14)+in_buf[600]*(5)+in_buf[601]*(0)+in_buf[602]*(17)+in_buf[603]*(22)+in_buf[604]*(6)+in_buf[605]*(0)+in_buf[606]*(-23)+in_buf[607]*(-29)+in_buf[608]*(-24)+in_buf[609]*(-21)+in_buf[610]*(-33)+in_buf[611]*(-49)+in_buf[612]*(-28)+in_buf[613]*(6)+in_buf[614]*(-6)+in_buf[615]*(2)+in_buf[616]*(0)+in_buf[617]*(9)+in_buf[618]*(-33)+in_buf[619]*(-21)+in_buf[620]*(-22)+in_buf[621]*(-1)+in_buf[622]*(25)+in_buf[623]*(2)+in_buf[624]*(-9)+in_buf[625]*(-8)+in_buf[626]*(3)+in_buf[627]*(6)+in_buf[628]*(0)+in_buf[629]*(-3)+in_buf[630]*(17)+in_buf[631]*(22)+in_buf[632]*(0)+in_buf[633]*(-17)+in_buf[634]*(-33)+in_buf[635]*(-45)+in_buf[636]*(-34)+in_buf[637]*(-7)+in_buf[638]*(-13)+in_buf[639]*(-38)+in_buf[640]*(-26)+in_buf[641]*(11)+in_buf[642]*(3)+in_buf[643]*(4)+in_buf[644]*(-1)+in_buf[645]*(2)+in_buf[646]*(-3)+in_buf[647]*(-24)+in_buf[648]*(-4)+in_buf[649]*(-16)+in_buf[650]*(-15)+in_buf[651]*(-18)+in_buf[652]*(-6)+in_buf[653]*(-1)+in_buf[654]*(1)+in_buf[655]*(-5)+in_buf[656]*(-5)+in_buf[657]*(2)+in_buf[658]*(13)+in_buf[659]*(7)+in_buf[660]*(-19)+in_buf[661]*(-29)+in_buf[662]*(-57)+in_buf[663]*(-47)+in_buf[664]*(-24)+in_buf[665]*(-25)+in_buf[666]*(-39)+in_buf[667]*(-22)+in_buf[668]*(-16)+in_buf[669]*(-15)+in_buf[670]*(19)+in_buf[671]*(-3)+in_buf[672]*(4)+in_buf[673]*(-2)+in_buf[674]*(11)+in_buf[675]*(11)+in_buf[676]*(-45)+in_buf[677]*(-24)+in_buf[678]*(-19)+in_buf[679]*(0)+in_buf[680]*(0)+in_buf[681]*(11)+in_buf[682]*(2)+in_buf[683]*(-22)+in_buf[684]*(0)+in_buf[685]*(-3)+in_buf[686]*(-15)+in_buf[687]*(-31)+in_buf[688]*(-27)+in_buf[689]*(-28)+in_buf[690]*(-59)+in_buf[691]*(-30)+in_buf[692]*(-25)+in_buf[693]*(-8)+in_buf[694]*(-29)+in_buf[695]*(-36)+in_buf[696]*(-9)+in_buf[697]*(14)+in_buf[698]*(18)+in_buf[699]*(-3)+in_buf[700]*(-1)+in_buf[701]*(-2)+in_buf[702]*(10)+in_buf[703]*(-17)+in_buf[704]*(-30)+in_buf[705]*(1)+in_buf[706]*(-1)+in_buf[707]*(12)+in_buf[708]*(19)+in_buf[709]*(28)+in_buf[710]*(9)+in_buf[711]*(-16)+in_buf[712]*(14)+in_buf[713]*(13)+in_buf[714]*(-13)+in_buf[715]*(-29)+in_buf[716]*(-16)+in_buf[717]*(-4)+in_buf[718]*(-37)+in_buf[719]*(-18)+in_buf[720]*(-16)+in_buf[721]*(-11)+in_buf[722]*(-8)+in_buf[723]*(-2)+in_buf[724]*(-2)+in_buf[725]*(0)+in_buf[726]*(3)+in_buf[727]*(2)+in_buf[728]*(-1)+in_buf[729]*(-1)+in_buf[730]*(1)+in_buf[731]*(-2)+in_buf[732]*(10)+in_buf[733]*(32)+in_buf[734]*(12)+in_buf[735]*(-25)+in_buf[736]*(-20)+in_buf[737]*(-20)+in_buf[738]*(4)+in_buf[739]*(8)+in_buf[740]*(-34)+in_buf[741]*(-67)+in_buf[742]*(-11)+in_buf[743]*(38)+in_buf[744]*(51)+in_buf[745]*(31)+in_buf[746]*(19)+in_buf[747]*(21)+in_buf[748]*(5)+in_buf[749]*(1)+in_buf[750]*(-15)+in_buf[751]*(-30)+in_buf[752]*(-3)+in_buf[753]*(-11)+in_buf[754]*(2)+in_buf[755]*(4)+in_buf[756]*(0)+in_buf[757]*(1)+in_buf[758]*(5)+in_buf[759]*(0)+in_buf[760]*(-9)+in_buf[761]*(-6)+in_buf[762]*(-6)+in_buf[763]*(1)+in_buf[764]*(5)+in_buf[765]*(-19)+in_buf[766]*(-9)+in_buf[767]*(-7)+in_buf[768]*(-15)+in_buf[769]*(-39)+in_buf[770]*(23)+in_buf[771]*(15)+in_buf[772]*(-5)+in_buf[773]*(6)+in_buf[774]*(20)+in_buf[775]*(9)+in_buf[776]*(1)+in_buf[777]*(-2)+in_buf[778]*(4)+in_buf[779]*(4)+in_buf[780]*(-1)+in_buf[781]*(4)+in_buf[782]*(0)+in_buf[783]*(-3);
assign in_buf_weight019=in_buf[0]*(4)+in_buf[1]*(-3)+in_buf[2]*(0)+in_buf[3]*(3)+in_buf[4]*(1)+in_buf[5]*(3)+in_buf[6]*(-4)+in_buf[7]*(1)+in_buf[8]*(-3)+in_buf[9]*(1)+in_buf[10]*(4)+in_buf[11]*(1)+in_buf[12]*(5)+in_buf[13]*(0)+in_buf[14]*(5)+in_buf[15]*(3)+in_buf[16]*(4)+in_buf[17]*(1)+in_buf[18]*(3)+in_buf[19]*(3)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(-2)+in_buf[23]*(-2)+in_buf[24]*(1)+in_buf[25]*(1)+in_buf[26]*(1)+in_buf[27]*(-1)+in_buf[28]*(0)+in_buf[29]*(-3)+in_buf[30]*(4)+in_buf[31]*(1)+in_buf[32]*(0)+in_buf[33]*(0)+in_buf[34]*(-9)+in_buf[35]*(-9)+in_buf[36]*(-10)+in_buf[37]*(-1)+in_buf[38]*(-3)+in_buf[39]*(9)+in_buf[40]*(8)+in_buf[41]*(24)+in_buf[42]*(23)+in_buf[43]*(0)+in_buf[44]*(4)+in_buf[45]*(8)+in_buf[46]*(2)+in_buf[47]*(-2)+in_buf[48]*(-12)+in_buf[49]*(-10)+in_buf[50]*(-6)+in_buf[51]*(-10)+in_buf[52]*(-3)+in_buf[53]*(-1)+in_buf[54]*(-2)+in_buf[55]*(1)+in_buf[56]*(-1)+in_buf[57]*(0)+in_buf[58]*(3)+in_buf[59]*(18)+in_buf[60]*(21)+in_buf[61]*(-9)+in_buf[62]*(-6)+in_buf[63]*(-3)+in_buf[64]*(-6)+in_buf[65]*(3)+in_buf[66]*(-3)+in_buf[67]*(-18)+in_buf[68]*(-37)+in_buf[69]*(-34)+in_buf[70]*(0)+in_buf[71]*(-9)+in_buf[72]*(-13)+in_buf[73]*(-22)+in_buf[74]*(-35)+in_buf[75]*(23)+in_buf[76]*(23)+in_buf[77]*(28)+in_buf[78]*(22)+in_buf[79]*(-5)+in_buf[80]*(0)+in_buf[81]*(-8)+in_buf[82]*(1)+in_buf[83]*(1)+in_buf[84]*(0)+in_buf[85]*(-3)+in_buf[86]*(7)+in_buf[87]*(13)+in_buf[88]*(-8)+in_buf[89]*(-16)+in_buf[90]*(-21)+in_buf[91]*(-6)+in_buf[92]*(-7)+in_buf[93]*(0)+in_buf[94]*(-3)+in_buf[95]*(-23)+in_buf[96]*(-40)+in_buf[97]*(-2)+in_buf[98]*(28)+in_buf[99]*(-1)+in_buf[100]*(-7)+in_buf[101]*(2)+in_buf[102]*(4)+in_buf[103]*(-5)+in_buf[104]*(-1)+in_buf[105]*(-13)+in_buf[106]*(-10)+in_buf[107]*(-9)+in_buf[108]*(-17)+in_buf[109]*(13)+in_buf[110]*(14)+in_buf[111]*(1)+in_buf[112]*(1)+in_buf[113]*(-4)+in_buf[114]*(-13)+in_buf[115]*(4)+in_buf[116]*(-20)+in_buf[117]*(-23)+in_buf[118]*(-32)+in_buf[119]*(-10)+in_buf[120]*(-15)+in_buf[121]*(-12)+in_buf[122]*(-19)+in_buf[123]*(-21)+in_buf[124]*(-12)+in_buf[125]*(-1)+in_buf[126]*(5)+in_buf[127]*(0)+in_buf[128]*(6)+in_buf[129]*(16)+in_buf[130]*(14)+in_buf[131]*(17)+in_buf[132]*(3)+in_buf[133]*(-1)+in_buf[134]*(-7)+in_buf[135]*(-2)+in_buf[136]*(0)+in_buf[137]*(3)+in_buf[138]*(-20)+in_buf[139]*(16)+in_buf[140]*(1)+in_buf[141]*(2)+in_buf[142]*(-14)+in_buf[143]*(10)+in_buf[144]*(-16)+in_buf[145]*(1)+in_buf[146]*(1)+in_buf[147]*(1)+in_buf[148]*(8)+in_buf[149]*(8)+in_buf[150]*(21)+in_buf[151]*(0)+in_buf[152]*(1)+in_buf[153]*(6)+in_buf[154]*(8)+in_buf[155]*(6)+in_buf[156]*(2)+in_buf[157]*(5)+in_buf[158]*(5)+in_buf[159]*(-3)+in_buf[160]*(-11)+in_buf[161]*(-3)+in_buf[162]*(2)+in_buf[163]*(-9)+in_buf[164]*(-1)+in_buf[165]*(16)+in_buf[166]*(-15)+in_buf[167]*(12)+in_buf[168]*(0)+in_buf[169]*(2)+in_buf[170]*(33)+in_buf[171]*(15)+in_buf[172]*(11)+in_buf[173]*(21)+in_buf[174]*(-6)+in_buf[175]*(4)+in_buf[176]*(-10)+in_buf[177]*(-15)+in_buf[178]*(10)+in_buf[179]*(26)+in_buf[180]*(33)+in_buf[181]*(17)+in_buf[182]*(-10)+in_buf[183]*(-16)+in_buf[184]*(-17)+in_buf[185]*(-7)+in_buf[186]*(-9)+in_buf[187]*(-3)+in_buf[188]*(-12)+in_buf[189]*(18)+in_buf[190]*(28)+in_buf[191]*(14)+in_buf[192]*(2)+in_buf[193]*(-22)+in_buf[194]*(-30)+in_buf[195]*(-11)+in_buf[196]*(1)+in_buf[197]*(5)+in_buf[198]*(27)+in_buf[199]*(12)+in_buf[200]*(-9)+in_buf[201]*(-7)+in_buf[202]*(-2)+in_buf[203]*(-14)+in_buf[204]*(-16)+in_buf[205]*(13)+in_buf[206]*(36)+in_buf[207]*(39)+in_buf[208]*(35)+in_buf[209]*(20)+in_buf[210]*(-6)+in_buf[211]*(-3)+in_buf[212]*(-9)+in_buf[213]*(9)+in_buf[214]*(19)+in_buf[215]*(5)+in_buf[216]*(0)+in_buf[217]*(15)+in_buf[218]*(28)+in_buf[219]*(26)+in_buf[220]*(18)+in_buf[221]*(17)+in_buf[222]*(4)+in_buf[223]*(-4)+in_buf[224]*(33)+in_buf[225]*(36)+in_buf[226]*(44)+in_buf[227]*(-30)+in_buf[228]*(-46)+in_buf[229]*(-25)+in_buf[230]*(0)+in_buf[231]*(-17)+in_buf[232]*(7)+in_buf[233]*(30)+in_buf[234]*(16)+in_buf[235]*(22)+in_buf[236]*(33)+in_buf[237]*(19)+in_buf[238]*(15)+in_buf[239]*(8)+in_buf[240]*(5)+in_buf[241]*(10)+in_buf[242]*(11)+in_buf[243]*(10)+in_buf[244]*(6)+in_buf[245]*(7)+in_buf[246]*(11)+in_buf[247]*(35)+in_buf[248]*(26)+in_buf[249]*(35)+in_buf[250]*(12)+in_buf[251]*(-13)+in_buf[252]*(16)+in_buf[253]*(30)+in_buf[254]*(6)+in_buf[255]*(-43)+in_buf[256]*(-54)+in_buf[257]*(-28)+in_buf[258]*(-17)+in_buf[259]*(0)+in_buf[260]*(-4)+in_buf[261]*(3)+in_buf[262]*(4)+in_buf[263]*(15)+in_buf[264]*(16)+in_buf[265]*(20)+in_buf[266]*(5)+in_buf[267]*(-19)+in_buf[268]*(-11)+in_buf[269]*(11)+in_buf[270]*(15)+in_buf[271]*(18)+in_buf[272]*(16)+in_buf[273]*(10)+in_buf[274]*(6)+in_buf[275]*(25)+in_buf[276]*(45)+in_buf[277]*(32)+in_buf[278]*(6)+in_buf[279]*(29)+in_buf[280]*(18)+in_buf[281]*(21)+in_buf[282]*(25)+in_buf[283]*(-25)+in_buf[284]*(-11)+in_buf[285]*(-10)+in_buf[286]*(-10)+in_buf[287]*(-4)+in_buf[288]*(-13)+in_buf[289]*(-2)+in_buf[290]*(4)+in_buf[291]*(14)+in_buf[292]*(4)+in_buf[293]*(7)+in_buf[294]*(-1)+in_buf[295]*(-8)+in_buf[296]*(-7)+in_buf[297]*(24)+in_buf[298]*(21)+in_buf[299]*(18)+in_buf[300]*(14)+in_buf[301]*(15)+in_buf[302]*(19)+in_buf[303]*(6)+in_buf[304]*(40)+in_buf[305]*(27)+in_buf[306]*(7)+in_buf[307]*(10)+in_buf[308]*(9)+in_buf[309]*(40)+in_buf[310]*(-27)+in_buf[311]*(-14)+in_buf[312]*(-24)+in_buf[313]*(-29)+in_buf[314]*(-1)+in_buf[315]*(14)+in_buf[316]*(-6)+in_buf[317]*(2)+in_buf[318]*(10)+in_buf[319]*(8)+in_buf[320]*(10)+in_buf[321]*(-5)+in_buf[322]*(-23)+in_buf[323]*(-25)+in_buf[324]*(-19)+in_buf[325]*(3)+in_buf[326]*(11)+in_buf[327]*(13)+in_buf[328]*(-1)+in_buf[329]*(12)+in_buf[330]*(13)+in_buf[331]*(5)+in_buf[332]*(9)+in_buf[333]*(7)+in_buf[334]*(-16)+in_buf[335]*(0)+in_buf[336]*(8)+in_buf[337]*(18)+in_buf[338]*(-11)+in_buf[339]*(-11)+in_buf[340]*(-38)+in_buf[341]*(-27)+in_buf[342]*(-7)+in_buf[343]*(-8)+in_buf[344]*(-6)+in_buf[345]*(10)+in_buf[346]*(17)+in_buf[347]*(24)+in_buf[348]*(23)+in_buf[349]*(-5)+in_buf[350]*(-35)+in_buf[351]*(-28)+in_buf[352]*(-19)+in_buf[353]*(-7)+in_buf[354]*(-2)+in_buf[355]*(-1)+in_buf[356]*(-6)+in_buf[357]*(-1)+in_buf[358]*(12)+in_buf[359]*(-24)+in_buf[360]*(-7)+in_buf[361]*(-20)+in_buf[362]*(-34)+in_buf[363]*(-23)+in_buf[364]*(3)+in_buf[365]*(25)+in_buf[366]*(49)+in_buf[367]*(3)+in_buf[368]*(-33)+in_buf[369]*(-19)+in_buf[370]*(8)+in_buf[371]*(10)+in_buf[372]*(5)+in_buf[373]*(20)+in_buf[374]*(19)+in_buf[375]*(15)+in_buf[376]*(7)+in_buf[377]*(-34)+in_buf[378]*(-15)+in_buf[379]*(-18)+in_buf[380]*(-16)+in_buf[381]*(1)+in_buf[382]*(5)+in_buf[383]*(-8)+in_buf[384]*(0)+in_buf[385]*(-3)+in_buf[386]*(3)+in_buf[387]*(0)+in_buf[388]*(8)+in_buf[389]*(-2)+in_buf[390]*(-29)+in_buf[391]*(-5)+in_buf[392]*(14)+in_buf[393]*(23)+in_buf[394]*(46)+in_buf[395]*(-5)+in_buf[396]*(-16)+in_buf[397]*(8)+in_buf[398]*(0)+in_buf[399]*(23)+in_buf[400]*(15)+in_buf[401]*(12)+in_buf[402]*(3)+in_buf[403]*(0)+in_buf[404]*(-9)+in_buf[405]*(-21)+in_buf[406]*(-13)+in_buf[407]*(-12)+in_buf[408]*(-18)+in_buf[409]*(7)+in_buf[410]*(-6)+in_buf[411]*(-4)+in_buf[412]*(-13)+in_buf[413]*(0)+in_buf[414]*(-3)+in_buf[415]*(2)+in_buf[416]*(23)+in_buf[417]*(23)+in_buf[418]*(-9)+in_buf[419]*(-2)+in_buf[420]*(12)+in_buf[421]*(-7)+in_buf[422]*(25)+in_buf[423]*(9)+in_buf[424]*(-15)+in_buf[425]*(-4)+in_buf[426]*(1)+in_buf[427]*(28)+in_buf[428]*(7)+in_buf[429]*(14)+in_buf[430]*(17)+in_buf[431]*(9)+in_buf[432]*(0)+in_buf[433]*(-14)+in_buf[434]*(-5)+in_buf[435]*(-7)+in_buf[436]*(-8)+in_buf[437]*(9)+in_buf[438]*(-7)+in_buf[439]*(-16)+in_buf[440]*(-7)+in_buf[441]*(7)+in_buf[442]*(11)+in_buf[443]*(6)+in_buf[444]*(14)+in_buf[445]*(5)+in_buf[446]*(1)+in_buf[447]*(9)+in_buf[448]*(13)+in_buf[449]*(-20)+in_buf[450]*(9)+in_buf[451]*(-10)+in_buf[452]*(-7)+in_buf[453]*(-6)+in_buf[454]*(7)+in_buf[455]*(23)+in_buf[456]*(23)+in_buf[457]*(17)+in_buf[458]*(16)+in_buf[459]*(3)+in_buf[460]*(-7)+in_buf[461]*(-4)+in_buf[462]*(3)+in_buf[463]*(-3)+in_buf[464]*(0)+in_buf[465]*(16)+in_buf[466]*(-9)+in_buf[467]*(-9)+in_buf[468]*(2)+in_buf[469]*(29)+in_buf[470]*(6)+in_buf[471]*(15)+in_buf[472]*(7)+in_buf[473]*(-8)+in_buf[474]*(2)+in_buf[475]*(14)+in_buf[476]*(3)+in_buf[477]*(-16)+in_buf[478]*(32)+in_buf[479]*(-29)+in_buf[480]*(11)+in_buf[481]*(12)+in_buf[482]*(15)+in_buf[483]*(14)+in_buf[484]*(23)+in_buf[485]*(26)+in_buf[486]*(5)+in_buf[487]*(-24)+in_buf[488]*(-14)+in_buf[489]*(6)+in_buf[490]*(11)+in_buf[491]*(-1)+in_buf[492]*(2)+in_buf[493]*(3)+in_buf[494]*(-3)+in_buf[495]*(-10)+in_buf[496]*(9)+in_buf[497]*(27)+in_buf[498]*(16)+in_buf[499]*(5)+in_buf[500]*(3)+in_buf[501]*(-19)+in_buf[502]*(-24)+in_buf[503]*(24)+in_buf[504]*(-13)+in_buf[505]*(-4)+in_buf[506]*(22)+in_buf[507]*(-24)+in_buf[508]*(7)+in_buf[509]*(22)+in_buf[510]*(15)+in_buf[511]*(20)+in_buf[512]*(18)+in_buf[513]*(4)+in_buf[514]*(-29)+in_buf[515]*(-42)+in_buf[516]*(-20)+in_buf[517]*(1)+in_buf[518]*(-4)+in_buf[519]*(-4)+in_buf[520]*(9)+in_buf[521]*(-4)+in_buf[522]*(1)+in_buf[523]*(-1)+in_buf[524]*(8)+in_buf[525]*(10)+in_buf[526]*(8)+in_buf[527]*(0)+in_buf[528]*(-8)+in_buf[529]*(-40)+in_buf[530]*(-12)+in_buf[531]*(7)+in_buf[532]*(-3)+in_buf[533]*(12)+in_buf[534]*(26)+in_buf[535]*(0)+in_buf[536]*(16)+in_buf[537]*(20)+in_buf[538]*(19)+in_buf[539]*(18)+in_buf[540]*(26)+in_buf[541]*(0)+in_buf[542]*(-38)+in_buf[543]*(-35)+in_buf[544]*(1)+in_buf[545]*(9)+in_buf[546]*(4)+in_buf[547]*(-1)+in_buf[548]*(-8)+in_buf[549]*(3)+in_buf[550]*(-7)+in_buf[551]*(0)+in_buf[552]*(4)+in_buf[553]*(18)+in_buf[554]*(8)+in_buf[555]*(-24)+in_buf[556]*(-30)+in_buf[557]*(-41)+in_buf[558]*(17)+in_buf[559]*(0)+in_buf[560]*(-1)+in_buf[561]*(13)+in_buf[562]*(29)+in_buf[563]*(24)+in_buf[564]*(8)+in_buf[565]*(13)+in_buf[566]*(10)+in_buf[567]*(15)+in_buf[568]*(29)+in_buf[569]*(10)+in_buf[570]*(-3)+in_buf[571]*(9)+in_buf[572]*(25)+in_buf[573]*(9)+in_buf[574]*(-16)+in_buf[575]*(-15)+in_buf[576]*(-16)+in_buf[577]*(-20)+in_buf[578]*(-24)+in_buf[579]*(-8)+in_buf[580]*(1)+in_buf[581]*(-2)+in_buf[582]*(-7)+in_buf[583]*(-41)+in_buf[584]*(-47)+in_buf[585]*(-51)+in_buf[586]*(22)+in_buf[587]*(0)+in_buf[588]*(-3)+in_buf[589]*(17)+in_buf[590]*(21)+in_buf[591]*(27)+in_buf[592]*(22)+in_buf[593]*(14)+in_buf[594]*(6)+in_buf[595]*(11)+in_buf[596]*(12)+in_buf[597]*(9)+in_buf[598]*(10)+in_buf[599]*(26)+in_buf[600]*(6)+in_buf[601]*(-10)+in_buf[602]*(-23)+in_buf[603]*(-19)+in_buf[604]*(-27)+in_buf[605]*(-28)+in_buf[606]*(-36)+in_buf[607]*(-20)+in_buf[608]*(-8)+in_buf[609]*(-17)+in_buf[610]*(4)+in_buf[611]*(-21)+in_buf[612]*(-37)+in_buf[613]*(-33)+in_buf[614]*(24)+in_buf[615]*(7)+in_buf[616]*(-6)+in_buf[617]*(2)+in_buf[618]*(24)+in_buf[619]*(32)+in_buf[620]*(0)+in_buf[621]*(-6)+in_buf[622]*(24)+in_buf[623]*(35)+in_buf[624]*(23)+in_buf[625]*(24)+in_buf[626]*(26)+in_buf[627]*(35)+in_buf[628]*(15)+in_buf[629]*(-8)+in_buf[630]*(-28)+in_buf[631]*(-15)+in_buf[632]*(-18)+in_buf[633]*(-31)+in_buf[634]*(-24)+in_buf[635]*(-7)+in_buf[636]*(-18)+in_buf[637]*(-14)+in_buf[638]*(3)+in_buf[639]*(-11)+in_buf[640]*(-27)+in_buf[641]*(-25)+in_buf[642]*(-4)+in_buf[643]*(2)+in_buf[644]*(2)+in_buf[645]*(0)+in_buf[646]*(-36)+in_buf[647]*(18)+in_buf[648]*(14)+in_buf[649]*(-10)+in_buf[650]*(36)+in_buf[651]*(42)+in_buf[652]*(27)+in_buf[653]*(20)+in_buf[654]*(27)+in_buf[655]*(26)+in_buf[656]*(13)+in_buf[657]*(-3)+in_buf[658]*(-9)+in_buf[659]*(-23)+in_buf[660]*(-21)+in_buf[661]*(-20)+in_buf[662]*(-34)+in_buf[663]*(-18)+in_buf[664]*(-32)+in_buf[665]*(-26)+in_buf[666]*(-22)+in_buf[667]*(-18)+in_buf[668]*(-30)+in_buf[669]*(-23)+in_buf[670]*(-19)+in_buf[671]*(-2)+in_buf[672]*(0)+in_buf[673]*(1)+in_buf[674]*(11)+in_buf[675]*(8)+in_buf[676]*(-6)+in_buf[677]*(13)+in_buf[678]*(22)+in_buf[679]*(12)+in_buf[680]*(0)+in_buf[681]*(9)+in_buf[682]*(1)+in_buf[683]*(17)+in_buf[684]*(10)+in_buf[685]*(12)+in_buf[686]*(-4)+in_buf[687]*(-21)+in_buf[688]*(-3)+in_buf[689]*(-7)+in_buf[690]*(-17)+in_buf[691]*(-40)+in_buf[692]*(-45)+in_buf[693]*(-17)+in_buf[694]*(-15)+in_buf[695]*(-30)+in_buf[696]*(-18)+in_buf[697]*(-4)+in_buf[698]*(-1)+in_buf[699]*(3)+in_buf[700]*(4)+in_buf[701]*(0)+in_buf[702]*(-36)+in_buf[703]*(24)+in_buf[704]*(16)+in_buf[705]*(-25)+in_buf[706]*(-4)+in_buf[707]*(-10)+in_buf[708]*(-19)+in_buf[709]*(-11)+in_buf[710]*(-4)+in_buf[711]*(2)+in_buf[712]*(-5)+in_buf[713]*(5)+in_buf[714]*(6)+in_buf[715]*(16)+in_buf[716]*(22)+in_buf[717]*(7)+in_buf[718]*(-12)+in_buf[719]*(-37)+in_buf[720]*(-36)+in_buf[721]*(-3)+in_buf[722]*(-10)+in_buf[723]*(-11)+in_buf[724]*(-26)+in_buf[725]*(8)+in_buf[726]*(13)+in_buf[727]*(0)+in_buf[728]*(-4)+in_buf[729]*(3)+in_buf[730]*(4)+in_buf[731]*(-12)+in_buf[732]*(-35)+in_buf[733]*(-55)+in_buf[734]*(-52)+in_buf[735]*(-23)+in_buf[736]*(3)+in_buf[737]*(-11)+in_buf[738]*(-11)+in_buf[739]*(3)+in_buf[740]*(16)+in_buf[741]*(12)+in_buf[742]*(-18)+in_buf[743]*(5)+in_buf[744]*(-2)+in_buf[745]*(-8)+in_buf[746]*(-18)+in_buf[747]*(3)+in_buf[748]*(-1)+in_buf[749]*(19)+in_buf[750]*(19)+in_buf[751]*(11)+in_buf[752]*(-24)+in_buf[753]*(14)+in_buf[754]*(-2)+in_buf[755]*(1)+in_buf[756]*(-1)+in_buf[757]*(0)+in_buf[758]*(4)+in_buf[759]*(3)+in_buf[760]*(33)+in_buf[761]*(27)+in_buf[762]*(4)+in_buf[763]*(-6)+in_buf[764]*(-13)+in_buf[765]*(-2)+in_buf[766]*(5)+in_buf[767]*(-9)+in_buf[768]*(-22)+in_buf[769]*(12)+in_buf[770]*(-24)+in_buf[771]*(-22)+in_buf[772]*(-6)+in_buf[773]*(-2)+in_buf[774]*(-7)+in_buf[775]*(-13)+in_buf[776]*(2)+in_buf[777]*(14)+in_buf[778]*(27)+in_buf[779]*(24)+in_buf[780]*(-3)+in_buf[781]*(-2)+in_buf[782]*(-2)+in_buf[783]*(0);
assign in_buf_weight020=in_buf[0]*(1)+in_buf[1]*(1)+in_buf[2]*(-2)+in_buf[3]*(3)+in_buf[4]*(1)+in_buf[5]*(1)+in_buf[6]*(2)+in_buf[7]*(-2)+in_buf[8]*(0)+in_buf[9]*(0)+in_buf[10]*(1)+in_buf[11]*(-1)+in_buf[12]*(-3)+in_buf[13]*(0)+in_buf[14]*(-1)+in_buf[15]*(4)+in_buf[16]*(4)+in_buf[17]*(2)+in_buf[18]*(4)+in_buf[19]*(3)+in_buf[20]*(-1)+in_buf[21]*(3)+in_buf[22]*(-1)+in_buf[23]*(-3)+in_buf[24]*(3)+in_buf[25]*(0)+in_buf[26]*(-1)+in_buf[27]*(-2)+in_buf[28]*(1)+in_buf[29]*(2)+in_buf[30]*(-3)+in_buf[31]*(0)+in_buf[32]*(0)+in_buf[33]*(-4)+in_buf[34]*(-6)+in_buf[35]*(-3)+in_buf[36]*(-2)+in_buf[37]*(-8)+in_buf[38]*(-6)+in_buf[39]*(-10)+in_buf[40]*(-14)+in_buf[41]*(-15)+in_buf[42]*(-2)+in_buf[43]*(-25)+in_buf[44]*(-24)+in_buf[45]*(-25)+in_buf[46]*(-10)+in_buf[47]*(-12)+in_buf[48]*(-16)+in_buf[49]*(-19)+in_buf[50]*(-14)+in_buf[51]*(-5)+in_buf[52]*(-2)+in_buf[53]*(1)+in_buf[54]*(2)+in_buf[55]*(-3)+in_buf[56]*(3)+in_buf[57]*(-2)+in_buf[58]*(-6)+in_buf[59]*(0)+in_buf[60]*(-1)+in_buf[61]*(-5)+in_buf[62]*(-8)+in_buf[63]*(-7)+in_buf[64]*(-12)+in_buf[65]*(-2)+in_buf[66]*(-2)+in_buf[67]*(3)+in_buf[68]*(-16)+in_buf[69]*(-43)+in_buf[70]*(-48)+in_buf[71]*(-24)+in_buf[72]*(-41)+in_buf[73]*(-18)+in_buf[74]*(-1)+in_buf[75]*(-25)+in_buf[76]*(-21)+in_buf[77]*(-11)+in_buf[78]*(-21)+in_buf[79]*(-19)+in_buf[80]*(-6)+in_buf[81]*(-7)+in_buf[82]*(4)+in_buf[83]*(0)+in_buf[84]*(-3)+in_buf[85]*(-2)+in_buf[86]*(2)+in_buf[87]*(-7)+in_buf[88]*(-2)+in_buf[89]*(0)+in_buf[90]*(-9)+in_buf[91]*(-9)+in_buf[92]*(-20)+in_buf[93]*(-20)+in_buf[94]*(-14)+in_buf[95]*(-9)+in_buf[96]*(-32)+in_buf[97]*(-60)+in_buf[98]*(-30)+in_buf[99]*(-29)+in_buf[100]*(-19)+in_buf[101]*(-12)+in_buf[102]*(-6)+in_buf[103]*(-19)+in_buf[104]*(-30)+in_buf[105]*(-13)+in_buf[106]*(-13)+in_buf[107]*(-20)+in_buf[108]*(0)+in_buf[109]*(-9)+in_buf[110]*(-4)+in_buf[111]*(4)+in_buf[112]*(3)+in_buf[113]*(2)+in_buf[114]*(0)+in_buf[115]*(-13)+in_buf[116]*(-14)+in_buf[117]*(-17)+in_buf[118]*(-13)+in_buf[119]*(-19)+in_buf[120]*(-32)+in_buf[121]*(-40)+in_buf[122]*(-30)+in_buf[123]*(16)+in_buf[124]*(-14)+in_buf[125]*(-25)+in_buf[126]*(-25)+in_buf[127]*(-27)+in_buf[128]*(-39)+in_buf[129]*(-43)+in_buf[130]*(-44)+in_buf[131]*(-52)+in_buf[132]*(-45)+in_buf[133]*(1)+in_buf[134]*(-11)+in_buf[135]*(-3)+in_buf[136]*(-13)+in_buf[137]*(-19)+in_buf[138]*(-14)+in_buf[139]*(-16)+in_buf[140]*(4)+in_buf[141]*(3)+in_buf[142]*(-14)+in_buf[143]*(-11)+in_buf[144]*(-29)+in_buf[145]*(-19)+in_buf[146]*(-31)+in_buf[147]*(-23)+in_buf[148]*(16)+in_buf[149]*(0)+in_buf[150]*(-3)+in_buf[151]*(12)+in_buf[152]*(3)+in_buf[153]*(-9)+in_buf[154]*(-12)+in_buf[155]*(-11)+in_buf[156]*(-42)+in_buf[157]*(-38)+in_buf[158]*(-30)+in_buf[159]*(-42)+in_buf[160]*(-40)+in_buf[161]*(-9)+in_buf[162]*(-2)+in_buf[163]*(30)+in_buf[164]*(18)+in_buf[165]*(-1)+in_buf[166]*(-30)+in_buf[167]*(-5)+in_buf[168]*(-2)+in_buf[169]*(-17)+in_buf[170]*(-2)+in_buf[171]*(-8)+in_buf[172]*(-10)+in_buf[173]*(-20)+in_buf[174]*(-8)+in_buf[175]*(10)+in_buf[176]*(12)+in_buf[177]*(10)+in_buf[178]*(-3)+in_buf[179]*(1)+in_buf[180]*(-3)+in_buf[181]*(10)+in_buf[182]*(4)+in_buf[183]*(1)+in_buf[184]*(14)+in_buf[185]*(15)+in_buf[186]*(-7)+in_buf[187]*(-25)+in_buf[188]*(-30)+in_buf[189]*(11)+in_buf[190]*(-2)+in_buf[191]*(-6)+in_buf[192]*(-9)+in_buf[193]*(-14)+in_buf[194]*(-16)+in_buf[195]*(-10)+in_buf[196]*(4)+in_buf[197]*(-35)+in_buf[198]*(-1)+in_buf[199]*(-10)+in_buf[200]*(-25)+in_buf[201]*(-21)+in_buf[202]*(8)+in_buf[203]*(-4)+in_buf[204]*(12)+in_buf[205]*(17)+in_buf[206]*(-1)+in_buf[207]*(-3)+in_buf[208]*(-1)+in_buf[209]*(10)+in_buf[210]*(6)+in_buf[211]*(7)+in_buf[212]*(13)+in_buf[213]*(11)+in_buf[214]*(-6)+in_buf[215]*(-14)+in_buf[216]*(-10)+in_buf[217]*(-7)+in_buf[218]*(-16)+in_buf[219]*(-10)+in_buf[220]*(2)+in_buf[221]*(-3)+in_buf[222]*(10)+in_buf[223]*(-6)+in_buf[224]*(-4)+in_buf[225]*(-13)+in_buf[226]*(-4)+in_buf[227]*(-13)+in_buf[228]*(-11)+in_buf[229]*(3)+in_buf[230]*(-9)+in_buf[231]*(-10)+in_buf[232]*(31)+in_buf[233]*(10)+in_buf[234]*(5)+in_buf[235]*(7)+in_buf[236]*(-13)+in_buf[237]*(-4)+in_buf[238]*(7)+in_buf[239]*(7)+in_buf[240]*(-7)+in_buf[241]*(-5)+in_buf[242]*(-6)+in_buf[243]*(-22)+in_buf[244]*(-26)+in_buf[245]*(-16)+in_buf[246]*(-23)+in_buf[247]*(-6)+in_buf[248]*(11)+in_buf[249]*(4)+in_buf[250]*(13)+in_buf[251]*(-4)+in_buf[252]*(6)+in_buf[253]*(7)+in_buf[254]*(26)+in_buf[255]*(17)+in_buf[256]*(-9)+in_buf[257]*(9)+in_buf[258]*(-7)+in_buf[259]*(1)+in_buf[260]*(6)+in_buf[261]*(3)+in_buf[262]*(7)+in_buf[263]*(0)+in_buf[264]*(4)+in_buf[265]*(0)+in_buf[266]*(2)+in_buf[267]*(13)+in_buf[268]*(-18)+in_buf[269]*(-9)+in_buf[270]*(-11)+in_buf[271]*(-24)+in_buf[272]*(-28)+in_buf[273]*(-8)+in_buf[274]*(-8)+in_buf[275]*(-12)+in_buf[276]*(6)+in_buf[277]*(-12)+in_buf[278]*(21)+in_buf[279]*(19)+in_buf[280]*(-1)+in_buf[281]*(-1)+in_buf[282]*(9)+in_buf[283]*(-16)+in_buf[284]*(-9)+in_buf[285]*(14)+in_buf[286]*(14)+in_buf[287]*(0)+in_buf[288]*(-2)+in_buf[289]*(1)+in_buf[290]*(-12)+in_buf[291]*(-1)+in_buf[292]*(10)+in_buf[293]*(2)+in_buf[294]*(15)+in_buf[295]*(16)+in_buf[296]*(2)+in_buf[297]*(-22)+in_buf[298]*(-27)+in_buf[299]*(-23)+in_buf[300]*(-4)+in_buf[301]*(10)+in_buf[302]*(8)+in_buf[303]*(-5)+in_buf[304]*(9)+in_buf[305]*(14)+in_buf[306]*(4)+in_buf[307]*(15)+in_buf[308]*(5)+in_buf[309]*(-13)+in_buf[310]*(-7)+in_buf[311]*(12)+in_buf[312]*(-11)+in_buf[313]*(6)+in_buf[314]*(2)+in_buf[315]*(11)+in_buf[316]*(10)+in_buf[317]*(-5)+in_buf[318]*(-9)+in_buf[319]*(3)+in_buf[320]*(21)+in_buf[321]*(1)+in_buf[322]*(5)+in_buf[323]*(26)+in_buf[324]*(17)+in_buf[325]*(7)+in_buf[326]*(-13)+in_buf[327]*(-2)+in_buf[328]*(1)+in_buf[329]*(4)+in_buf[330]*(11)+in_buf[331]*(-3)+in_buf[332]*(-5)+in_buf[333]*(-10)+in_buf[334]*(-47)+in_buf[335]*(27)+in_buf[336]*(7)+in_buf[337]*(-6)+in_buf[338]*(8)+in_buf[339]*(19)+in_buf[340]*(3)+in_buf[341]*(3)+in_buf[342]*(6)+in_buf[343]*(16)+in_buf[344]*(7)+in_buf[345]*(1)+in_buf[346]*(-3)+in_buf[347]*(8)+in_buf[348]*(9)+in_buf[349]*(0)+in_buf[350]*(18)+in_buf[351]*(43)+in_buf[352]*(28)+in_buf[353]*(18)+in_buf[354]*(13)+in_buf[355]*(4)+in_buf[356]*(9)+in_buf[357]*(3)+in_buf[358]*(-4)+in_buf[359]*(-20)+in_buf[360]*(-33)+in_buf[361]*(-16)+in_buf[362]*(-9)+in_buf[363]*(25)+in_buf[364]*(-25)+in_buf[365]*(4)+in_buf[366]*(16)+in_buf[367]*(19)+in_buf[368]*(26)+in_buf[369]*(1)+in_buf[370]*(24)+in_buf[371]*(19)+in_buf[372]*(6)+in_buf[373]*(0)+in_buf[374]*(13)+in_buf[375]*(2)+in_buf[376]*(15)+in_buf[377]*(15)+in_buf[378]*(21)+in_buf[379]*(27)+in_buf[380]*(31)+in_buf[381]*(13)+in_buf[382]*(15)+in_buf[383]*(16)+in_buf[384]*(13)+in_buf[385]*(1)+in_buf[386]*(-17)+in_buf[387]*(-32)+in_buf[388]*(-27)+in_buf[389]*(-14)+in_buf[390]*(-12)+in_buf[391]*(-1)+in_buf[392]*(-14)+in_buf[393]*(7)+in_buf[394]*(4)+in_buf[395]*(13)+in_buf[396]*(26)+in_buf[397]*(-5)+in_buf[398]*(4)+in_buf[399]*(13)+in_buf[400]*(2)+in_buf[401]*(3)+in_buf[402]*(14)+in_buf[403]*(13)+in_buf[404]*(23)+in_buf[405]*(18)+in_buf[406]*(12)+in_buf[407]*(16)+in_buf[408]*(18)+in_buf[409]*(16)+in_buf[410]*(26)+in_buf[411]*(16)+in_buf[412]*(8)+in_buf[413]*(-23)+in_buf[414]*(-16)+in_buf[415]*(-22)+in_buf[416]*(-23)+in_buf[417]*(-6)+in_buf[418]*(-29)+in_buf[419]*(13)+in_buf[420]*(-8)+in_buf[421]*(-1)+in_buf[422]*(-24)+in_buf[423]*(24)+in_buf[424]*(24)+in_buf[425]*(-2)+in_buf[426]*(-31)+in_buf[427]*(-23)+in_buf[428]*(-7)+in_buf[429]*(0)+in_buf[430]*(28)+in_buf[431]*(28)+in_buf[432]*(16)+in_buf[433]*(14)+in_buf[434]*(6)+in_buf[435]*(24)+in_buf[436]*(21)+in_buf[437]*(38)+in_buf[438]*(20)+in_buf[439]*(12)+in_buf[440]*(-5)+in_buf[441]*(-8)+in_buf[442]*(-4)+in_buf[443]*(1)+in_buf[444]*(16)+in_buf[445]*(8)+in_buf[446]*(7)+in_buf[447]*(-15)+in_buf[448]*(8)+in_buf[449]*(-2)+in_buf[450]*(-8)+in_buf[451]*(12)+in_buf[452]*(26)+in_buf[453]*(2)+in_buf[454]*(-20)+in_buf[455]*(-15)+in_buf[456]*(3)+in_buf[457]*(-4)+in_buf[458]*(20)+in_buf[459]*(28)+in_buf[460]*(10)+in_buf[461]*(-3)+in_buf[462]*(5)+in_buf[463]*(32)+in_buf[464]*(30)+in_buf[465]*(22)+in_buf[466]*(-2)+in_buf[467]*(-6)+in_buf[468]*(-11)+in_buf[469]*(-11)+in_buf[470]*(-4)+in_buf[471]*(8)+in_buf[472]*(3)+in_buf[473]*(5)+in_buf[474]*(8)+in_buf[475]*(-10)+in_buf[476]*(-1)+in_buf[477]*(-6)+in_buf[478]*(8)+in_buf[479]*(-4)+in_buf[480]*(8)+in_buf[481]*(14)+in_buf[482]*(-5)+in_buf[483]*(-26)+in_buf[484]*(-13)+in_buf[485]*(-9)+in_buf[486]*(2)+in_buf[487]*(-9)+in_buf[488]*(-12)+in_buf[489]*(0)+in_buf[490]*(11)+in_buf[491]*(23)+in_buf[492]*(13)+in_buf[493]*(-8)+in_buf[494]*(-10)+in_buf[495]*(-24)+in_buf[496]*(-22)+in_buf[497]*(-13)+in_buf[498]*(-13)+in_buf[499]*(20)+in_buf[500]*(1)+in_buf[501]*(35)+in_buf[502]*(-1)+in_buf[503]*(-16)+in_buf[504]*(1)+in_buf[505]*(-2)+in_buf[506]*(10)+in_buf[507]*(-8)+in_buf[508]*(-6)+in_buf[509]*(-2)+in_buf[510]*(-17)+in_buf[511]*(-32)+in_buf[512]*(-24)+in_buf[513]*(-35)+in_buf[514]*(-24)+in_buf[515]*(-20)+in_buf[516]*(-30)+in_buf[517]*(0)+in_buf[518]*(9)+in_buf[519]*(4)+in_buf[520]*(-10)+in_buf[521]*(-33)+in_buf[522]*(-35)+in_buf[523]*(-44)+in_buf[524]*(-38)+in_buf[525]*(-23)+in_buf[526]*(-19)+in_buf[527]*(-7)+in_buf[528]*(-24)+in_buf[529]*(14)+in_buf[530]*(27)+in_buf[531]*(2)+in_buf[532]*(-11)+in_buf[533]*(-11)+in_buf[534]*(0)+in_buf[535]*(-34)+in_buf[536]*(-27)+in_buf[537]*(-21)+in_buf[538]*(-14)+in_buf[539]*(-14)+in_buf[540]*(-27)+in_buf[541]*(-41)+in_buf[542]*(-41)+in_buf[543]*(-32)+in_buf[544]*(-24)+in_buf[545]*(2)+in_buf[546]*(6)+in_buf[547]*(0)+in_buf[548]*(-12)+in_buf[549]*(-31)+in_buf[550]*(-53)+in_buf[551]*(-44)+in_buf[552]*(-39)+in_buf[553]*(-10)+in_buf[554]*(-24)+in_buf[555]*(-32)+in_buf[556]*(-51)+in_buf[557]*(-12)+in_buf[558]*(-2)+in_buf[559]*(4)+in_buf[560]*(-2)+in_buf[561]*(-3)+in_buf[562]*(-14)+in_buf[563]*(-46)+in_buf[564]*(-22)+in_buf[565]*(-13)+in_buf[566]*(-14)+in_buf[567]*(-30)+in_buf[568]*(-24)+in_buf[569]*(-27)+in_buf[570]*(-11)+in_buf[571]*(-15)+in_buf[572]*(-13)+in_buf[573]*(2)+in_buf[574]*(1)+in_buf[575]*(-15)+in_buf[576]*(-7)+in_buf[577]*(-38)+in_buf[578]*(-42)+in_buf[579]*(-44)+in_buf[580]*(-33)+in_buf[581]*(-16)+in_buf[582]*(-17)+in_buf[583]*(-25)+in_buf[584]*(-6)+in_buf[585]*(0)+in_buf[586]*(0)+in_buf[587]*(-4)+in_buf[588]*(13)+in_buf[589]*(-1)+in_buf[590]*(-14)+in_buf[591]*(-37)+in_buf[592]*(-15)+in_buf[593]*(0)+in_buf[594]*(-26)+in_buf[595]*(-25)+in_buf[596]*(0)+in_buf[597]*(17)+in_buf[598]*(8)+in_buf[599]*(1)+in_buf[600]*(2)+in_buf[601]*(-5)+in_buf[602]*(-17)+in_buf[603]*(-21)+in_buf[604]*(-25)+in_buf[605]*(-38)+in_buf[606]*(-33)+in_buf[607]*(-32)+in_buf[608]*(-22)+in_buf[609]*(-10)+in_buf[610]*(-21)+in_buf[611]*(-17)+in_buf[612]*(-5)+in_buf[613]*(-20)+in_buf[614]*(-13)+in_buf[615]*(1)+in_buf[616]*(11)+in_buf[617]*(7)+in_buf[618]*(-12)+in_buf[619]*(-6)+in_buf[620]*(-15)+in_buf[621]*(-31)+in_buf[622]*(-30)+in_buf[623]*(-26)+in_buf[624]*(12)+in_buf[625]*(2)+in_buf[626]*(12)+in_buf[627]*(0)+in_buf[628]*(3)+in_buf[629]*(-3)+in_buf[630]*(2)+in_buf[631]*(-15)+in_buf[632]*(-16)+in_buf[633]*(-13)+in_buf[634]*(-12)+in_buf[635]*(-25)+in_buf[636]*(-11)+in_buf[637]*(-27)+in_buf[638]*(-20)+in_buf[639]*(-11)+in_buf[640]*(-8)+in_buf[641]*(6)+in_buf[642]*(-21)+in_buf[643]*(1)+in_buf[644]*(-1)+in_buf[645]*(4)+in_buf[646]*(-23)+in_buf[647]*(4)+in_buf[648]*(-34)+in_buf[649]*(-48)+in_buf[650]*(-39)+in_buf[651]*(-24)+in_buf[652]*(0)+in_buf[653]*(-11)+in_buf[654]*(-4)+in_buf[655]*(-4)+in_buf[656]*(9)+in_buf[657]*(13)+in_buf[658]*(7)+in_buf[659]*(-12)+in_buf[660]*(1)+in_buf[661]*(8)+in_buf[662]*(10)+in_buf[663]*(-5)+in_buf[664]*(5)+in_buf[665]*(1)+in_buf[666]*(-9)+in_buf[667]*(-1)+in_buf[668]*(10)+in_buf[669]*(-4)+in_buf[670]*(2)+in_buf[671]*(-3)+in_buf[672]*(4)+in_buf[673]*(-2)+in_buf[674]*(-20)+in_buf[675]*(-18)+in_buf[676]*(-15)+in_buf[677]*(-20)+in_buf[678]*(-28)+in_buf[679]*(-20)+in_buf[680]*(3)+in_buf[681]*(-12)+in_buf[682]*(-13)+in_buf[683]*(-9)+in_buf[684]*(-24)+in_buf[685]*(1)+in_buf[686]*(-6)+in_buf[687]*(-9)+in_buf[688]*(-10)+in_buf[689]*(17)+in_buf[690]*(19)+in_buf[691]*(8)+in_buf[692]*(15)+in_buf[693]*(4)+in_buf[694]*(0)+in_buf[695]*(18)+in_buf[696]*(3)+in_buf[697]*(12)+in_buf[698]*(5)+in_buf[699]*(-2)+in_buf[700]*(-1)+in_buf[701]*(-3)+in_buf[702]*(3)+in_buf[703]*(-6)+in_buf[704]*(-8)+in_buf[705]*(9)+in_buf[706]*(-7)+in_buf[707]*(-7)+in_buf[708]*(6)+in_buf[709]*(-6)+in_buf[710]*(-17)+in_buf[711]*(-5)+in_buf[712]*(-15)+in_buf[713]*(-18)+in_buf[714]*(-1)+in_buf[715]*(-12)+in_buf[716]*(-12)+in_buf[717]*(9)+in_buf[718]*(5)+in_buf[719]*(-15)+in_buf[720]*(-15)+in_buf[721]*(-20)+in_buf[722]*(-21)+in_buf[723]*(-11)+in_buf[724]*(-15)+in_buf[725]*(16)+in_buf[726]*(5)+in_buf[727]*(2)+in_buf[728]*(-1)+in_buf[729]*(-1)+in_buf[730]*(0)+in_buf[731]*(10)+in_buf[732]*(17)+in_buf[733]*(18)+in_buf[734]*(16)+in_buf[735]*(12)+in_buf[736]*(11)+in_buf[737]*(17)+in_buf[738]*(32)+in_buf[739]*(12)+in_buf[740]*(9)+in_buf[741]*(9)+in_buf[742]*(33)+in_buf[743]*(7)+in_buf[744]*(10)+in_buf[745]*(12)+in_buf[746]*(9)+in_buf[747]*(8)+in_buf[748]*(11)+in_buf[749]*(0)+in_buf[750]*(-6)+in_buf[751]*(-13)+in_buf[752]*(-2)+in_buf[753]*(0)+in_buf[754]*(-3)+in_buf[755]*(0)+in_buf[756]*(-1)+in_buf[757]*(0)+in_buf[758]*(1)+in_buf[759]*(2)+in_buf[760]*(1)+in_buf[761]*(11)+in_buf[762]*(16)+in_buf[763]*(12)+in_buf[764]*(9)+in_buf[765]*(12)+in_buf[766]*(39)+in_buf[767]*(22)+in_buf[768]*(14)+in_buf[769]*(12)+in_buf[770]*(57)+in_buf[771]*(24)+in_buf[772]*(20)+in_buf[773]*(32)+in_buf[774]*(28)+in_buf[775]*(39)+in_buf[776]*(23)+in_buf[777]*(11)+in_buf[778]*(14)+in_buf[779]*(0)+in_buf[780]*(3)+in_buf[781]*(-1)+in_buf[782]*(4)+in_buf[783]*(4);
assign in_buf_weight021=in_buf[0]*(1)+in_buf[1]*(3)+in_buf[2]*(1)+in_buf[3]*(1)+in_buf[4]*(-3)+in_buf[5]*(-1)+in_buf[6]*(1)+in_buf[7]*(-3)+in_buf[8]*(1)+in_buf[9]*(2)+in_buf[10]*(4)+in_buf[11]*(3)+in_buf[12]*(0)+in_buf[13]*(-3)+in_buf[14]*(1)+in_buf[15]*(0)+in_buf[16]*(0)+in_buf[17]*(3)+in_buf[18]*(4)+in_buf[19]*(0)+in_buf[20]*(0)+in_buf[21]*(-2)+in_buf[22]*(4)+in_buf[23]*(0)+in_buf[24]*(0)+in_buf[25]*(3)+in_buf[26]*(-1)+in_buf[27]*(4)+in_buf[28]*(2)+in_buf[29]*(2)+in_buf[30]*(4)+in_buf[31]*(-3)+in_buf[32]*(0)+in_buf[33]*(-2)+in_buf[34]*(-2)+in_buf[35]*(2)+in_buf[36]*(-2)+in_buf[37]*(-2)+in_buf[38]*(-7)+in_buf[39]*(-3)+in_buf[40]*(-7)+in_buf[41]*(-10)+in_buf[42]*(-2)+in_buf[43]*(0)+in_buf[44]*(9)+in_buf[45]*(1)+in_buf[46]*(-3)+in_buf[47]*(-8)+in_buf[48]*(-9)+in_buf[49]*(-5)+in_buf[50]*(-2)+in_buf[51]*(-4)+in_buf[52]*(-2)+in_buf[53]*(0)+in_buf[54]*(-2)+in_buf[55]*(-1)+in_buf[56]*(-3)+in_buf[57]*(-4)+in_buf[58]*(-3)+in_buf[59]*(2)+in_buf[60]*(2)+in_buf[61]*(-2)+in_buf[62]*(1)+in_buf[63]*(-6)+in_buf[64]*(16)+in_buf[65]*(20)+in_buf[66]*(3)+in_buf[67]*(-16)+in_buf[68]*(-9)+in_buf[69]*(-6)+in_buf[70]*(-16)+in_buf[71]*(-17)+in_buf[72]*(-29)+in_buf[73]*(-30)+in_buf[74]*(-11)+in_buf[75]*(-6)+in_buf[76]*(4)+in_buf[77]*(5)+in_buf[78]*(-3)+in_buf[79]*(-9)+in_buf[80]*(0)+in_buf[81]*(-1)+in_buf[82]*(4)+in_buf[83]*(3)+in_buf[84]*(2)+in_buf[85]*(1)+in_buf[86]*(8)+in_buf[87]*(0)+in_buf[88]*(-2)+in_buf[89]*(0)+in_buf[90]*(5)+in_buf[91]*(9)+in_buf[92]*(-4)+in_buf[93]*(17)+in_buf[94]*(6)+in_buf[95]*(-18)+in_buf[96]*(-20)+in_buf[97]*(-6)+in_buf[98]*(27)+in_buf[99]*(17)+in_buf[100]*(23)+in_buf[101]*(10)+in_buf[102]*(8)+in_buf[103]*(14)+in_buf[104]*(-18)+in_buf[105]*(-16)+in_buf[106]*(-20)+in_buf[107]*(-35)+in_buf[108]*(-18)+in_buf[109]*(5)+in_buf[110]*(6)+in_buf[111]*(1)+in_buf[112]*(1)+in_buf[113]*(0)+in_buf[114]*(8)+in_buf[115]*(-24)+in_buf[116]*(-8)+in_buf[117]*(19)+in_buf[118]*(65)+in_buf[119]*(49)+in_buf[120]*(25)+in_buf[121]*(30)+in_buf[122]*(9)+in_buf[123]*(15)+in_buf[124]*(0)+in_buf[125]*(-3)+in_buf[126]*(-7)+in_buf[127]*(-12)+in_buf[128]*(-6)+in_buf[129]*(7)+in_buf[130]*(1)+in_buf[131]*(5)+in_buf[132]*(-3)+in_buf[133]*(-1)+in_buf[134]*(4)+in_buf[135]*(0)+in_buf[136]*(4)+in_buf[137]*(22)+in_buf[138]*(28)+in_buf[139]*(15)+in_buf[140]*(-3)+in_buf[141]*(0)+in_buf[142]*(8)+in_buf[143]*(17)+in_buf[144]*(-5)+in_buf[145]*(-1)+in_buf[146]*(16)+in_buf[147]*(12)+in_buf[148]*(15)+in_buf[149]*(11)+in_buf[150]*(26)+in_buf[151]*(28)+in_buf[152]*(25)+in_buf[153]*(16)+in_buf[154]*(-7)+in_buf[155]*(-17)+in_buf[156]*(0)+in_buf[157]*(-1)+in_buf[158]*(-4)+in_buf[159]*(-6)+in_buf[160]*(4)+in_buf[161]*(6)+in_buf[162]*(21)+in_buf[163]*(27)+in_buf[164]*(15)+in_buf[165]*(19)+in_buf[166]*(17)+in_buf[167]*(10)+in_buf[168]*(-3)+in_buf[169]*(4)+in_buf[170]*(19)+in_buf[171]*(8)+in_buf[172]*(-2)+in_buf[173]*(-11)+in_buf[174]*(3)+in_buf[175]*(4)+in_buf[176]*(-12)+in_buf[177]*(2)+in_buf[178]*(25)+in_buf[179]*(8)+in_buf[180]*(13)+in_buf[181]*(13)+in_buf[182]*(11)+in_buf[183]*(-1)+in_buf[184]*(-3)+in_buf[185]*(-10)+in_buf[186]*(8)+in_buf[187]*(10)+in_buf[188]*(3)+in_buf[189]*(18)+in_buf[190]*(25)+in_buf[191]*(32)+in_buf[192]*(35)+in_buf[193]*(8)+in_buf[194]*(-14)+in_buf[195]*(14)+in_buf[196]*(-3)+in_buf[197]*(21)+in_buf[198]*(13)+in_buf[199]*(20)+in_buf[200]*(11)+in_buf[201]*(24)+in_buf[202]*(1)+in_buf[203]*(15)+in_buf[204]*(8)+in_buf[205]*(0)+in_buf[206]*(-4)+in_buf[207]*(5)+in_buf[208]*(3)+in_buf[209]*(8)+in_buf[210]*(26)+in_buf[211]*(12)+in_buf[212]*(6)+in_buf[213]*(6)+in_buf[214]*(16)+in_buf[215]*(24)+in_buf[216]*(17)+in_buf[217]*(21)+in_buf[218]*(16)+in_buf[219]*(28)+in_buf[220]*(23)+in_buf[221]*(0)+in_buf[222]*(-16)+in_buf[223]*(7)+in_buf[224]*(0)+in_buf[225]*(14)+in_buf[226]*(-11)+in_buf[227]*(-20)+in_buf[228]*(29)+in_buf[229]*(16)+in_buf[230]*(4)+in_buf[231]*(-2)+in_buf[232]*(1)+in_buf[233]*(0)+in_buf[234]*(-17)+in_buf[235]*(-14)+in_buf[236]*(-16)+in_buf[237]*(-11)+in_buf[238]*(19)+in_buf[239]*(12)+in_buf[240]*(5)+in_buf[241]*(13)+in_buf[242]*(26)+in_buf[243]*(18)+in_buf[244]*(9)+in_buf[245]*(19)+in_buf[246]*(19)+in_buf[247]*(31)+in_buf[248]*(21)+in_buf[249]*(3)+in_buf[250]*(1)+in_buf[251]*(-4)+in_buf[252]*(-3)+in_buf[253]*(14)+in_buf[254]*(-5)+in_buf[255]*(-13)+in_buf[256]*(24)+in_buf[257]*(19)+in_buf[258]*(-7)+in_buf[259]*(-3)+in_buf[260]*(-12)+in_buf[261]*(-4)+in_buf[262]*(-17)+in_buf[263]*(-20)+in_buf[264]*(-11)+in_buf[265]*(-19)+in_buf[266]*(-5)+in_buf[267]*(-13)+in_buf[268]*(-11)+in_buf[269]*(-9)+in_buf[270]*(4)+in_buf[271]*(-8)+in_buf[272]*(-3)+in_buf[273]*(10)+in_buf[274]*(17)+in_buf[275]*(21)+in_buf[276]*(26)+in_buf[277]*(30)+in_buf[278]*(-6)+in_buf[279]*(11)+in_buf[280]*(-3)+in_buf[281]*(4)+in_buf[282]*(-1)+in_buf[283]*(9)+in_buf[284]*(-2)+in_buf[285]*(0)+in_buf[286]*(-17)+in_buf[287]*(-4)+in_buf[288]*(3)+in_buf[289]*(-4)+in_buf[290]*(-10)+in_buf[291]*(-13)+in_buf[292]*(-1)+in_buf[293]*(-12)+in_buf[294]*(-14)+in_buf[295]*(-22)+in_buf[296]*(-10)+in_buf[297]*(-14)+in_buf[298]*(-15)+in_buf[299]*(-29)+in_buf[300]*(-7)+in_buf[301]*(15)+in_buf[302]*(11)+in_buf[303]*(-10)+in_buf[304]*(6)+in_buf[305]*(17)+in_buf[306]*(35)+in_buf[307]*(10)+in_buf[308]*(-3)+in_buf[309]*(16)+in_buf[310]*(-10)+in_buf[311]*(-18)+in_buf[312]*(-8)+in_buf[313]*(-18)+in_buf[314]*(-18)+in_buf[315]*(-13)+in_buf[316]*(5)+in_buf[317]*(-25)+in_buf[318]*(-17)+in_buf[319]*(-16)+in_buf[320]*(-37)+in_buf[321]*(-37)+in_buf[322]*(-33)+in_buf[323]*(-25)+in_buf[324]*(-19)+in_buf[325]*(-22)+in_buf[326]*(-21)+in_buf[327]*(-24)+in_buf[328]*(-6)+in_buf[329]*(14)+in_buf[330]*(5)+in_buf[331]*(-2)+in_buf[332]*(-8)+in_buf[333]*(-6)+in_buf[334]*(18)+in_buf[335]*(19)+in_buf[336]*(0)+in_buf[337]*(10)+in_buf[338]*(0)+in_buf[339]*(-27)+in_buf[340]*(-5)+in_buf[341]*(-11)+in_buf[342]*(-7)+in_buf[343]*(-24)+in_buf[344]*(-12)+in_buf[345]*(-17)+in_buf[346]*(-16)+in_buf[347]*(-24)+in_buf[348]*(-32)+in_buf[349]*(-26)+in_buf[350]*(-12)+in_buf[351]*(-18)+in_buf[352]*(-33)+in_buf[353]*(-28)+in_buf[354]*(-29)+in_buf[355]*(-18)+in_buf[356]*(7)+in_buf[357]*(14)+in_buf[358]*(-7)+in_buf[359]*(9)+in_buf[360]*(-14)+in_buf[361]*(-11)+in_buf[362]*(-1)+in_buf[363]*(-1)+in_buf[364]*(0)+in_buf[365]*(1)+in_buf[366]*(0)+in_buf[367]*(4)+in_buf[368]*(23)+in_buf[369]*(-3)+in_buf[370]*(3)+in_buf[371]*(-5)+in_buf[372]*(0)+in_buf[373]*(-6)+in_buf[374]*(-11)+in_buf[375]*(-23)+in_buf[376]*(-24)+in_buf[377]*(1)+in_buf[378]*(3)+in_buf[379]*(-12)+in_buf[380]*(-24)+in_buf[381]*(-43)+in_buf[382]*(-28)+in_buf[383]*(-3)+in_buf[384]*(3)+in_buf[385]*(25)+in_buf[386]*(4)+in_buf[387]*(-3)+in_buf[388]*(-11)+in_buf[389]*(7)+in_buf[390]*(13)+in_buf[391]*(1)+in_buf[392]*(10)+in_buf[393]*(-3)+in_buf[394]*(-6)+in_buf[395]*(11)+in_buf[396]*(27)+in_buf[397]*(4)+in_buf[398]*(3)+in_buf[399]*(19)+in_buf[400]*(16)+in_buf[401]*(4)+in_buf[402]*(-5)+in_buf[403]*(-5)+in_buf[404]*(-8)+in_buf[405]*(19)+in_buf[406]*(27)+in_buf[407]*(3)+in_buf[408]*(-29)+in_buf[409]*(-50)+in_buf[410]*(-21)+in_buf[411]*(-11)+in_buf[412]*(9)+in_buf[413]*(22)+in_buf[414]*(2)+in_buf[415]*(-4)+in_buf[416]*(-7)+in_buf[417]*(-9)+in_buf[418]*(33)+in_buf[419]*(14)+in_buf[420]*(3)+in_buf[421]*(-8)+in_buf[422]*(-8)+in_buf[423]*(33)+in_buf[424]*(10)+in_buf[425]*(0)+in_buf[426]*(2)+in_buf[427]*(8)+in_buf[428]*(15)+in_buf[429]*(11)+in_buf[430]*(3)+in_buf[431]*(-9)+in_buf[432]*(6)+in_buf[433]*(22)+in_buf[434]*(27)+in_buf[435]*(-2)+in_buf[436]*(-34)+in_buf[437]*(-44)+in_buf[438]*(-24)+in_buf[439]*(0)+in_buf[440]*(15)+in_buf[441]*(27)+in_buf[442]*(-1)+in_buf[443]*(-4)+in_buf[444]*(8)+in_buf[445]*(-12)+in_buf[446]*(34)+in_buf[447]*(27)+in_buf[448]*(-4)+in_buf[449]*(-8)+in_buf[450]*(-4)+in_buf[451]*(26)+in_buf[452]*(8)+in_buf[453]*(19)+in_buf[454]*(0)+in_buf[455]*(3)+in_buf[456]*(-3)+in_buf[457]*(-4)+in_buf[458]*(3)+in_buf[459]*(-3)+in_buf[460]*(4)+in_buf[461]*(24)+in_buf[462]*(6)+in_buf[463]*(-14)+in_buf[464]*(-34)+in_buf[465]*(-44)+in_buf[466]*(-20)+in_buf[467]*(17)+in_buf[468]*(19)+in_buf[469]*(10)+in_buf[470]*(0)+in_buf[471]*(4)+in_buf[472]*(9)+in_buf[473]*(0)+in_buf[474]*(47)+in_buf[475]*(29)+in_buf[476]*(2)+in_buf[477]*(-8)+in_buf[478]*(-5)+in_buf[479]*(34)+in_buf[480]*(17)+in_buf[481]*(8)+in_buf[482]*(10)+in_buf[483]*(2)+in_buf[484]*(-18)+in_buf[485]*(-13)+in_buf[486]*(-11)+in_buf[487]*(-17)+in_buf[488]*(-4)+in_buf[489]*(-1)+in_buf[490]*(-21)+in_buf[491]*(-53)+in_buf[492]*(-52)+in_buf[493]*(-30)+in_buf[494]*(0)+in_buf[495]*(16)+in_buf[496]*(11)+in_buf[497]*(0)+in_buf[498]*(0)+in_buf[499]*(-11)+in_buf[500]*(-5)+in_buf[501]*(28)+in_buf[502]*(28)+in_buf[503]*(24)+in_buf[504]*(4)+in_buf[505]*(-9)+in_buf[506]*(-15)+in_buf[507]*(27)+in_buf[508]*(4)+in_buf[509]*(-1)+in_buf[510]*(8)+in_buf[511]*(17)+in_buf[512]*(5)+in_buf[513]*(-2)+in_buf[514]*(-23)+in_buf[515]*(-29)+in_buf[516]*(-7)+in_buf[517]*(-23)+in_buf[518]*(-43)+in_buf[519]*(-55)+in_buf[520]*(-21)+in_buf[521]*(-11)+in_buf[522]*(12)+in_buf[523]*(11)+in_buf[524]*(6)+in_buf[525]*(5)+in_buf[526]*(0)+in_buf[527]*(-7)+in_buf[528]*(-3)+in_buf[529]*(24)+in_buf[530]*(15)+in_buf[531]*(32)+in_buf[532]*(-11)+in_buf[533]*(0)+in_buf[534]*(7)+in_buf[535]*(8)+in_buf[536]*(-16)+in_buf[537]*(0)+in_buf[538]*(16)+in_buf[539]*(16)+in_buf[540]*(4)+in_buf[541]*(-1)+in_buf[542]*(-9)+in_buf[543]*(4)+in_buf[544]*(4)+in_buf[545]*(-3)+in_buf[546]*(-24)+in_buf[547]*(-29)+in_buf[548]*(-8)+in_buf[549]*(5)+in_buf[550]*(4)+in_buf[551]*(-7)+in_buf[552]*(6)+in_buf[553]*(1)+in_buf[554]*(-10)+in_buf[555]*(-29)+in_buf[556]*(-14)+in_buf[557]*(12)+in_buf[558]*(44)+in_buf[559]*(30)+in_buf[560]*(1)+in_buf[561]*(3)+in_buf[562]*(12)+in_buf[563]*(34)+in_buf[564]*(-20)+in_buf[565]*(20)+in_buf[566]*(9)+in_buf[567]*(9)+in_buf[568]*(7)+in_buf[569]*(14)+in_buf[570]*(3)+in_buf[571]*(23)+in_buf[572]*(14)+in_buf[573]*(13)+in_buf[574]*(11)+in_buf[575]*(12)+in_buf[576]*(21)+in_buf[577]*(1)+in_buf[578]*(-5)+in_buf[579]*(-1)+in_buf[580]*(-9)+in_buf[581]*(-7)+in_buf[582]*(-3)+in_buf[583]*(-4)+in_buf[584]*(-20)+in_buf[585]*(-5)+in_buf[586]*(33)+in_buf[587]*(-12)+in_buf[588]*(0)+in_buf[589]*(15)+in_buf[590]*(10)+in_buf[591]*(37)+in_buf[592]*(-6)+in_buf[593]*(-12)+in_buf[594]*(-9)+in_buf[595]*(0)+in_buf[596]*(6)+in_buf[597]*(7)+in_buf[598]*(12)+in_buf[599]*(20)+in_buf[600]*(23)+in_buf[601]*(35)+in_buf[602]*(45)+in_buf[603]*(39)+in_buf[604]*(24)+in_buf[605]*(5)+in_buf[606]*(1)+in_buf[607]*(-3)+in_buf[608]*(-3)+in_buf[609]*(-1)+in_buf[610]*(13)+in_buf[611]*(23)+in_buf[612]*(5)+in_buf[613]*(15)+in_buf[614]*(18)+in_buf[615]*(2)+in_buf[616]*(0)+in_buf[617]*(2)+in_buf[618]*(8)+in_buf[619]*(45)+in_buf[620]*(-4)+in_buf[621]*(-14)+in_buf[622]*(-6)+in_buf[623]*(0)+in_buf[624]*(18)+in_buf[625]*(20)+in_buf[626]*(12)+in_buf[627]*(20)+in_buf[628]*(17)+in_buf[629]*(31)+in_buf[630]*(35)+in_buf[631]*(24)+in_buf[632]*(23)+in_buf[633]*(19)+in_buf[634]*(19)+in_buf[635]*(19)+in_buf[636]*(4)+in_buf[637]*(9)+in_buf[638]*(25)+in_buf[639]*(17)+in_buf[640]*(8)+in_buf[641]*(6)+in_buf[642]*(-10)+in_buf[643]*(8)+in_buf[644]*(-2)+in_buf[645]*(-1)+in_buf[646]*(3)+in_buf[647]*(33)+in_buf[648]*(1)+in_buf[649]*(21)+in_buf[650]*(6)+in_buf[651]*(-10)+in_buf[652]*(-4)+in_buf[653]*(10)+in_buf[654]*(13)+in_buf[655]*(22)+in_buf[656]*(20)+in_buf[657]*(14)+in_buf[658]*(24)+in_buf[659]*(27)+in_buf[660]*(15)+in_buf[661]*(22)+in_buf[662]*(14)+in_buf[663]*(17)+in_buf[664]*(13)+in_buf[665]*(10)+in_buf[666]*(25)+in_buf[667]*(5)+in_buf[668]*(1)+in_buf[669]*(11)+in_buf[670]*(-4)+in_buf[671]*(-3)+in_buf[672]*(3)+in_buf[673]*(2)+in_buf[674]*(-7)+in_buf[675]*(2)+in_buf[676]*(0)+in_buf[677]*(-5)+in_buf[678]*(11)+in_buf[679]*(15)+in_buf[680]*(5)+in_buf[681]*(16)+in_buf[682]*(13)+in_buf[683]*(9)+in_buf[684]*(15)+in_buf[685]*(19)+in_buf[686]*(24)+in_buf[687]*(29)+in_buf[688]*(0)+in_buf[689]*(9)+in_buf[690]*(15)+in_buf[691]*(-7)+in_buf[692]*(1)+in_buf[693]*(23)+in_buf[694]*(16)+in_buf[695]*(0)+in_buf[696]*(22)+in_buf[697]*(21)+in_buf[698]*(9)+in_buf[699]*(-1)+in_buf[700]*(-1)+in_buf[701]*(1)+in_buf[702]*(1)+in_buf[703]*(1)+in_buf[704]*(-16)+in_buf[705]*(-15)+in_buf[706]*(-7)+in_buf[707]*(0)+in_buf[708]*(5)+in_buf[709]*(7)+in_buf[710]*(19)+in_buf[711]*(7)+in_buf[712]*(2)+in_buf[713]*(-23)+in_buf[714]*(-18)+in_buf[715]*(3)+in_buf[716]*(1)+in_buf[717]*(-7)+in_buf[718]*(-6)+in_buf[719]*(0)+in_buf[720]*(0)+in_buf[721]*(11)+in_buf[722]*(20)+in_buf[723]*(1)+in_buf[724]*(11)+in_buf[725]*(8)+in_buf[726]*(5)+in_buf[727]*(2)+in_buf[728]*(0)+in_buf[729]*(-1)+in_buf[730]*(0)+in_buf[731]*(3)+in_buf[732]*(-1)+in_buf[733]*(1)+in_buf[734]*(8)+in_buf[735]*(0)+in_buf[736]*(-2)+in_buf[737]*(-9)+in_buf[738]*(3)+in_buf[739]*(11)+in_buf[740]*(37)+in_buf[741]*(18)+in_buf[742]*(-15)+in_buf[743]*(-5)+in_buf[744]*(-12)+in_buf[745]*(-30)+in_buf[746]*(-22)+in_buf[747]*(0)+in_buf[748]*(-23)+in_buf[749]*(-19)+in_buf[750]*(-9)+in_buf[751]*(-8)+in_buf[752]*(0)+in_buf[753]*(-3)+in_buf[754]*(1)+in_buf[755]*(-2)+in_buf[756]*(4)+in_buf[757]*(-1)+in_buf[758]*(3)+in_buf[759]*(2)+in_buf[760]*(0)+in_buf[761]*(2)+in_buf[762]*(-6)+in_buf[763]*(0)+in_buf[764]*(-3)+in_buf[765]*(2)+in_buf[766]*(-5)+in_buf[767]*(-7)+in_buf[768]*(-1)+in_buf[769]*(-14)+in_buf[770]*(-11)+in_buf[771]*(-6)+in_buf[772]*(-8)+in_buf[773]*(-4)+in_buf[774]*(-3)+in_buf[775]*(0)+in_buf[776]*(1)+in_buf[777]*(-8)+in_buf[778]*(-11)+in_buf[779]*(-7)+in_buf[780]*(4)+in_buf[781]*(3)+in_buf[782]*(0)+in_buf[783]*(1);
assign in_buf_weight022=in_buf[0]*(0)+in_buf[1]*(-3)+in_buf[2]*(0)+in_buf[3]*(2)+in_buf[4]*(-3)+in_buf[5]*(-2)+in_buf[6]*(3)+in_buf[7]*(-3)+in_buf[8]*(-1)+in_buf[9]*(-2)+in_buf[10]*(0)+in_buf[11]*(2)+in_buf[12]*(1)+in_buf[13]*(-5)+in_buf[14]*(-5)+in_buf[15]*(-2)+in_buf[16]*(-1)+in_buf[17]*(1)+in_buf[18]*(3)+in_buf[19]*(3)+in_buf[20]*(0)+in_buf[21]*(1)+in_buf[22]*(4)+in_buf[23]*(-1)+in_buf[24]*(2)+in_buf[25]*(-3)+in_buf[26]*(3)+in_buf[27]*(-2)+in_buf[28]*(-1)+in_buf[29]*(0)+in_buf[30]*(1)+in_buf[31]*(-1)+in_buf[32]*(-3)+in_buf[33]*(-1)+in_buf[34]*(-3)+in_buf[35]*(-1)+in_buf[36]*(-1)+in_buf[37]*(-5)+in_buf[38]*(-8)+in_buf[39]*(-28)+in_buf[40]*(-31)+in_buf[41]*(-24)+in_buf[42]*(-5)+in_buf[43]*(-26)+in_buf[44]*(-31)+in_buf[45]*(-28)+in_buf[46]*(-18)+in_buf[47]*(-25)+in_buf[48]*(-21)+in_buf[49]*(-15)+in_buf[50]*(-16)+in_buf[51]*(-8)+in_buf[52]*(0)+in_buf[53]*(-1)+in_buf[54]*(4)+in_buf[55]*(0)+in_buf[56]*(1)+in_buf[57]*(-3)+in_buf[58]*(-5)+in_buf[59]*(-19)+in_buf[60]*(-25)+in_buf[61]*(0)+in_buf[62]*(-8)+in_buf[63]*(-5)+in_buf[64]*(-6)+in_buf[65]*(-16)+in_buf[66]*(-12)+in_buf[67]*(-6)+in_buf[68]*(-8)+in_buf[69]*(-19)+in_buf[70]*(-20)+in_buf[71]*(-43)+in_buf[72]*(-41)+in_buf[73]*(-14)+in_buf[74]*(-52)+in_buf[75]*(-52)+in_buf[76]*(-42)+in_buf[77]*(-40)+in_buf[78]*(-37)+in_buf[79]*(-29)+in_buf[80]*(-17)+in_buf[81]*(-2)+in_buf[82]*(-2)+in_buf[83]*(-1)+in_buf[84]*(3)+in_buf[85]*(3)+in_buf[86]*(17)+in_buf[87]*(-23)+in_buf[88]*(-27)+in_buf[89]*(-34)+in_buf[90]*(-19)+in_buf[91]*(-10)+in_buf[92]*(-34)+in_buf[93]*(-39)+in_buf[94]*(-27)+in_buf[95]*(-30)+in_buf[96]*(-31)+in_buf[97]*(-50)+in_buf[98]*(-43)+in_buf[99]*(-81)+in_buf[100]*(-40)+in_buf[101]*(18)+in_buf[102]*(7)+in_buf[103]*(7)+in_buf[104]*(-15)+in_buf[105]*(-47)+in_buf[106]*(-25)+in_buf[107]*(-30)+in_buf[108]*(-32)+in_buf[109]*(-29)+in_buf[110]*(-20)+in_buf[111]*(-1)+in_buf[112]*(-1)+in_buf[113]*(0)+in_buf[114]*(14)+in_buf[115]*(19)+in_buf[116]*(-24)+in_buf[117]*(-22)+in_buf[118]*(2)+in_buf[119]*(-19)+in_buf[120]*(-38)+in_buf[121]*(-56)+in_buf[122]*(-58)+in_buf[123]*(-30)+in_buf[124]*(-35)+in_buf[125]*(-27)+in_buf[126]*(-62)+in_buf[127]*(-36)+in_buf[128]*(-17)+in_buf[129]*(-28)+in_buf[130]*(-20)+in_buf[131]*(-2)+in_buf[132]*(-13)+in_buf[133]*(-5)+in_buf[134]*(-3)+in_buf[135]*(-22)+in_buf[136]*(-33)+in_buf[137]*(-48)+in_buf[138]*(-15)+in_buf[139]*(-26)+in_buf[140]*(-3)+in_buf[141]*(4)+in_buf[142]*(-15)+in_buf[143]*(1)+in_buf[144]*(-33)+in_buf[145]*(-6)+in_buf[146]*(17)+in_buf[147]*(9)+in_buf[148]*(10)+in_buf[149]*(4)+in_buf[150]*(-5)+in_buf[151]*(0)+in_buf[152]*(-7)+in_buf[153]*(-22)+in_buf[154]*(-25)+in_buf[155]*(-19)+in_buf[156]*(-10)+in_buf[157]*(-9)+in_buf[158]*(-4)+in_buf[159]*(-15)+in_buf[160]*(-21)+in_buf[161]*(-13)+in_buf[162]*(-7)+in_buf[163]*(-15)+in_buf[164]*(-10)+in_buf[165]*(-13)+in_buf[166]*(-45)+in_buf[167]*(-10)+in_buf[168]*(2)+in_buf[169]*(-22)+in_buf[170]*(-15)+in_buf[171]*(14)+in_buf[172]*(-21)+in_buf[173]*(12)+in_buf[174]*(18)+in_buf[175]*(6)+in_buf[176]*(-11)+in_buf[177]*(10)+in_buf[178]*(-6)+in_buf[179]*(-3)+in_buf[180]*(-5)+in_buf[181]*(-12)+in_buf[182]*(3)+in_buf[183]*(3)+in_buf[184]*(10)+in_buf[185]*(28)+in_buf[186]*(19)+in_buf[187]*(9)+in_buf[188]*(16)+in_buf[189]*(4)+in_buf[190]*(-9)+in_buf[191]*(-4)+in_buf[192]*(-3)+in_buf[193]*(-18)+in_buf[194]*(-16)+in_buf[195]*(-26)+in_buf[196]*(4)+in_buf[197]*(-19)+in_buf[198]*(-8)+in_buf[199]*(36)+in_buf[200]*(-20)+in_buf[201]*(-22)+in_buf[202]*(-12)+in_buf[203]*(-18)+in_buf[204]*(-19)+in_buf[205]*(0)+in_buf[206]*(0)+in_buf[207]*(-10)+in_buf[208]*(-9)+in_buf[209]*(3)+in_buf[210]*(9)+in_buf[211]*(11)+in_buf[212]*(14)+in_buf[213]*(19)+in_buf[214]*(7)+in_buf[215]*(18)+in_buf[216]*(23)+in_buf[217]*(12)+in_buf[218]*(-6)+in_buf[219]*(14)+in_buf[220]*(12)+in_buf[221]*(-20)+in_buf[222]*(-8)+in_buf[223]*(-23)+in_buf[224]*(-34)+in_buf[225]*(10)+in_buf[226]*(-13)+in_buf[227]*(20)+in_buf[228]*(-7)+in_buf[229]*(-6)+in_buf[230]*(-8)+in_buf[231]*(-12)+in_buf[232]*(8)+in_buf[233]*(13)+in_buf[234]*(4)+in_buf[235]*(-9)+in_buf[236]*(-7)+in_buf[237]*(5)+in_buf[238]*(7)+in_buf[239]*(15)+in_buf[240]*(2)+in_buf[241]*(12)+in_buf[242]*(9)+in_buf[243]*(-3)+in_buf[244]*(-3)+in_buf[245]*(-1)+in_buf[246]*(-11)+in_buf[247]*(-8)+in_buf[248]*(23)+in_buf[249]*(8)+in_buf[250]*(10)+in_buf[251]*(-3)+in_buf[252]*(16)+in_buf[253]*(27)+in_buf[254]*(-3)+in_buf[255]*(-14)+in_buf[256]*(-15)+in_buf[257]*(-15)+in_buf[258]*(-10)+in_buf[259]*(-9)+in_buf[260]*(14)+in_buf[261]*(10)+in_buf[262]*(18)+in_buf[263]*(-2)+in_buf[264]*(1)+in_buf[265]*(0)+in_buf[266]*(4)+in_buf[267]*(26)+in_buf[268]*(6)+in_buf[269]*(8)+in_buf[270]*(7)+in_buf[271]*(-5)+in_buf[272]*(0)+in_buf[273]*(-6)+in_buf[274]*(-7)+in_buf[275]*(-15)+in_buf[276]*(-3)+in_buf[277]*(-17)+in_buf[278]*(22)+in_buf[279]*(23)+in_buf[280]*(10)+in_buf[281]*(12)+in_buf[282]*(-13)+in_buf[283]*(-38)+in_buf[284]*(-13)+in_buf[285]*(-5)+in_buf[286]*(-24)+in_buf[287]*(-33)+in_buf[288]*(-6)+in_buf[289]*(25)+in_buf[290]*(7)+in_buf[291]*(5)+in_buf[292]*(0)+in_buf[293]*(-21)+in_buf[294]*(0)+in_buf[295]*(23)+in_buf[296]*(17)+in_buf[297]*(-3)+in_buf[298]*(-5)+in_buf[299]*(8)+in_buf[300]*(2)+in_buf[301]*(-11)+in_buf[302]*(-17)+in_buf[303]*(-15)+in_buf[304]*(0)+in_buf[305]*(28)+in_buf[306]*(-10)+in_buf[307]*(20)+in_buf[308]*(14)+in_buf[309]*(-36)+in_buf[310]*(27)+in_buf[311]*(5)+in_buf[312]*(-4)+in_buf[313]*(3)+in_buf[314]*(-22)+in_buf[315]*(-14)+in_buf[316]*(19)+in_buf[317]*(25)+in_buf[318]*(15)+in_buf[319]*(4)+in_buf[320]*(-18)+in_buf[321]*(-27)+in_buf[322]*(11)+in_buf[323]*(24)+in_buf[324]*(28)+in_buf[325]*(11)+in_buf[326]*(10)+in_buf[327]*(7)+in_buf[328]*(-2)+in_buf[329]*(-7)+in_buf[330]*(-9)+in_buf[331]*(-18)+in_buf[332]*(13)+in_buf[333]*(-3)+in_buf[334]*(-54)+in_buf[335]*(31)+in_buf[336]*(11)+in_buf[337]*(-11)+in_buf[338]*(43)+in_buf[339]*(17)+in_buf[340]*(0)+in_buf[341]*(-7)+in_buf[342]*(0)+in_buf[343]*(0)+in_buf[344]*(10)+in_buf[345]*(0)+in_buf[346]*(3)+in_buf[347]*(-13)+in_buf[348]*(-37)+in_buf[349]*(-20)+in_buf[350]*(22)+in_buf[351]*(36)+in_buf[352]*(26)+in_buf[353]*(10)+in_buf[354]*(15)+in_buf[355]*(15)+in_buf[356]*(-1)+in_buf[357]*(-2)+in_buf[358]*(-15)+in_buf[359]*(-6)+in_buf[360]*(-16)+in_buf[361]*(0)+in_buf[362]*(-13)+in_buf[363]*(40)+in_buf[364]*(-18)+in_buf[365]*(-8)+in_buf[366]*(25)+in_buf[367]*(21)+in_buf[368]*(34)+in_buf[369]*(-25)+in_buf[370]*(-6)+in_buf[371]*(30)+in_buf[372]*(9)+in_buf[373]*(0)+in_buf[374]*(0)+in_buf[375]*(-23)+in_buf[376]*(-32)+in_buf[377]*(-7)+in_buf[378]*(27)+in_buf[379]*(34)+in_buf[380]*(14)+in_buf[381]*(3)+in_buf[382]*(8)+in_buf[383]*(5)+in_buf[384]*(8)+in_buf[385]*(3)+in_buf[386]*(-10)+in_buf[387]*(-33)+in_buf[388]*(-29)+in_buf[389]*(-20)+in_buf[390]*(-48)+in_buf[391]*(-22)+in_buf[392]*(-5)+in_buf[393]*(-14)+in_buf[394]*(-2)+in_buf[395]*(23)+in_buf[396]*(30)+in_buf[397]*(-31)+in_buf[398]*(-6)+in_buf[399]*(26)+in_buf[400]*(18)+in_buf[401]*(-1)+in_buf[402]*(-10)+in_buf[403]*(-16)+in_buf[404]*(-13)+in_buf[405]*(13)+in_buf[406]*(31)+in_buf[407]*(24)+in_buf[408]*(23)+in_buf[409]*(15)+in_buf[410]*(14)+in_buf[411]*(19)+in_buf[412]*(14)+in_buf[413]*(-18)+in_buf[414]*(-20)+in_buf[415]*(-25)+in_buf[416]*(-36)+in_buf[417]*(-31)+in_buf[418]*(-40)+in_buf[419]*(-10)+in_buf[420]*(-1)+in_buf[421]*(1)+in_buf[422]*(-13)+in_buf[423]*(-12)+in_buf[424]*(10)+in_buf[425]*(-2)+in_buf[426]*(1)+in_buf[427]*(26)+in_buf[428]*(24)+in_buf[429]*(7)+in_buf[430]*(22)+in_buf[431]*(13)+in_buf[432]*(0)+in_buf[433]*(5)+in_buf[434]*(18)+in_buf[435]*(29)+in_buf[436]*(22)+in_buf[437]*(29)+in_buf[438]*(16)+in_buf[439]*(1)+in_buf[440]*(-2)+in_buf[441]*(-1)+in_buf[442]*(1)+in_buf[443]*(-6)+in_buf[444]*(-21)+in_buf[445]*(-33)+in_buf[446]*(-17)+in_buf[447]*(-16)+in_buf[448]*(11)+in_buf[449]*(-1)+in_buf[450]*(-23)+in_buf[451]*(-47)+in_buf[452]*(-5)+in_buf[453]*(0)+in_buf[454]*(14)+in_buf[455]*(31)+in_buf[456]*(43)+in_buf[457]*(20)+in_buf[458]*(15)+in_buf[459]*(11)+in_buf[460]*(10)+in_buf[461]*(14)+in_buf[462]*(14)+in_buf[463]*(14)+in_buf[464]*(24)+in_buf[465]*(11)+in_buf[466]*(-7)+in_buf[467]*(-14)+in_buf[468]*(-8)+in_buf[469]*(-6)+in_buf[470]*(-2)+in_buf[471]*(11)+in_buf[472]*(-11)+in_buf[473]*(-32)+in_buf[474]*(-41)+in_buf[475]*(-35)+in_buf[476]*(1)+in_buf[477]*(-6)+in_buf[478]*(-39)+in_buf[479]*(-19)+in_buf[480]*(-21)+in_buf[481]*(-12)+in_buf[482]*(9)+in_buf[483]*(29)+in_buf[484]*(35)+in_buf[485]*(31)+in_buf[486]*(22)+in_buf[487]*(19)+in_buf[488]*(25)+in_buf[489]*(20)+in_buf[490]*(18)+in_buf[491]*(7)+in_buf[492]*(5)+in_buf[493]*(-10)+in_buf[494]*(-8)+in_buf[495]*(-16)+in_buf[496]*(-2)+in_buf[497]*(3)+in_buf[498]*(7)+in_buf[499]*(2)+in_buf[500]*(-6)+in_buf[501]*(5)+in_buf[502]*(-27)+in_buf[503]*(-31)+in_buf[504]*(36)+in_buf[505]*(1)+in_buf[506]*(-27)+in_buf[507]*(-15)+in_buf[508]*(-28)+in_buf[509]*(-24)+in_buf[510]*(-27)+in_buf[511]*(5)+in_buf[512]*(8)+in_buf[513]*(2)+in_buf[514]*(6)+in_buf[515]*(23)+in_buf[516]*(4)+in_buf[517]*(24)+in_buf[518]*(5)+in_buf[519]*(-11)+in_buf[520]*(-21)+in_buf[521]*(-17)+in_buf[522]*(-27)+in_buf[523]*(-26)+in_buf[524]*(-17)+in_buf[525]*(1)+in_buf[526]*(-4)+in_buf[527]*(-20)+in_buf[528]*(-39)+in_buf[529]*(1)+in_buf[530]*(22)+in_buf[531]*(17)+in_buf[532]*(12)+in_buf[533]*(-19)+in_buf[534]*(-3)+in_buf[535]*(-44)+in_buf[536]*(-46)+in_buf[537]*(-43)+in_buf[538]*(-28)+in_buf[539]*(-4)+in_buf[540]*(-11)+in_buf[541]*(-21)+in_buf[542]*(-10)+in_buf[543]*(-3)+in_buf[544]*(1)+in_buf[545]*(14)+in_buf[546]*(0)+in_buf[547]*(-13)+in_buf[548]*(-26)+in_buf[549]*(-36)+in_buf[550]*(-48)+in_buf[551]*(-30)+in_buf[552]*(-37)+in_buf[553]*(-6)+in_buf[554]*(-15)+in_buf[555]*(-36)+in_buf[556]*(-50)+in_buf[557]*(3)+in_buf[558]*(-31)+in_buf[559]*(16)+in_buf[560]*(0)+in_buf[561]*(-26)+in_buf[562]*(-34)+in_buf[563]*(-55)+in_buf[564]*(-42)+in_buf[565]*(-23)+in_buf[566]*(-35)+in_buf[567]*(-43)+in_buf[568]*(-39)+in_buf[569]*(-32)+in_buf[570]*(-25)+in_buf[571]*(-14)+in_buf[572]*(-6)+in_buf[573]*(7)+in_buf[574]*(3)+in_buf[575]*(-11)+in_buf[576]*(-11)+in_buf[577]*(-28)+in_buf[578]*(-25)+in_buf[579]*(-31)+in_buf[580]*(-36)+in_buf[581]*(-8)+in_buf[582]*(6)+in_buf[583]*(-11)+in_buf[584]*(-4)+in_buf[585]*(11)+in_buf[586]*(-35)+in_buf[587]*(4)+in_buf[588]*(19)+in_buf[589]*(7)+in_buf[590]*(-28)+in_buf[591]*(-23)+in_buf[592]*(-9)+in_buf[593]*(-8)+in_buf[594]*(-27)+in_buf[595]*(-33)+in_buf[596]*(-20)+in_buf[597]*(-5)+in_buf[598]*(-3)+in_buf[599]*(-24)+in_buf[600]*(-15)+in_buf[601]*(-4)+in_buf[602]*(-3)+in_buf[603]*(-8)+in_buf[604]*(-19)+in_buf[605]*(-30)+in_buf[606]*(-29)+in_buf[607]*(-42)+in_buf[608]*(-20)+in_buf[609]*(16)+in_buf[610]*(2)+in_buf[611]*(-9)+in_buf[612]*(4)+in_buf[613]*(-7)+in_buf[614]*(-32)+in_buf[615]*(0)+in_buf[616]*(20)+in_buf[617]*(17)+in_buf[618]*(-16)+in_buf[619]*(-9)+in_buf[620]*(13)+in_buf[621]*(15)+in_buf[622]*(-1)+in_buf[623]*(-1)+in_buf[624]*(2)+in_buf[625]*(-4)+in_buf[626]*(3)+in_buf[627]*(-16)+in_buf[628]*(-17)+in_buf[629]*(-7)+in_buf[630]*(8)+in_buf[631]*(-8)+in_buf[632]*(-24)+in_buf[633]*(-23)+in_buf[634]*(-32)+in_buf[635]*(-37)+in_buf[636]*(-9)+in_buf[637]*(12)+in_buf[638]*(-10)+in_buf[639]*(-5)+in_buf[640]*(-2)+in_buf[641]*(3)+in_buf[642]*(-33)+in_buf[643]*(2)+in_buf[644]*(-2)+in_buf[645]*(4)+in_buf[646]*(-30)+in_buf[647]*(-30)+in_buf[648]*(-19)+in_buf[649]*(8)+in_buf[650]*(17)+in_buf[651]*(11)+in_buf[652]*(15)+in_buf[653]*(2)+in_buf[654]*(-1)+in_buf[655]*(-5)+in_buf[656]*(-8)+in_buf[657]*(-3)+in_buf[658]*(0)+in_buf[659]*(-15)+in_buf[660]*(-12)+in_buf[661]*(-5)+in_buf[662]*(-16)+in_buf[663]*(-31)+in_buf[664]*(-7)+in_buf[665]*(1)+in_buf[666]*(14)+in_buf[667]*(10)+in_buf[668]*(8)+in_buf[669]*(-8)+in_buf[670]*(8)+in_buf[671]*(4)+in_buf[672]*(0)+in_buf[673]*(-1)+in_buf[674]*(-12)+in_buf[675]*(-35)+in_buf[676]*(14)+in_buf[677]*(14)+in_buf[678]*(6)+in_buf[679]*(18)+in_buf[680]*(19)+in_buf[681]*(-2)+in_buf[682]*(-10)+in_buf[683]*(-2)+in_buf[684]*(-18)+in_buf[685]*(-3)+in_buf[686]*(-13)+in_buf[687]*(-5)+in_buf[688]*(-12)+in_buf[689]*(-21)+in_buf[690]*(-31)+in_buf[691]*(-45)+in_buf[692]*(-35)+in_buf[693]*(-3)+in_buf[694]*(9)+in_buf[695]*(37)+in_buf[696]*(-7)+in_buf[697]*(15)+in_buf[698]*(4)+in_buf[699]*(-1)+in_buf[700]*(0)+in_buf[701]*(1)+in_buf[702]*(19)+in_buf[703]*(22)+in_buf[704]*(13)+in_buf[705]*(24)+in_buf[706]*(-8)+in_buf[707]*(-9)+in_buf[708]*(9)+in_buf[709]*(4)+in_buf[710]*(-12)+in_buf[711]*(-2)+in_buf[712]*(-8)+in_buf[713]*(-17)+in_buf[714]*(1)+in_buf[715]*(-8)+in_buf[716]*(-6)+in_buf[717]*(-28)+in_buf[718]*(-37)+in_buf[719]*(-34)+in_buf[720]*(-25)+in_buf[721]*(-18)+in_buf[722]*(-14)+in_buf[723]*(5)+in_buf[724]*(-7)+in_buf[725]*(5)+in_buf[726]*(-5)+in_buf[727]*(-2)+in_buf[728]*(0)+in_buf[729]*(-3)+in_buf[730]*(1)+in_buf[731]*(14)+in_buf[732]*(9)+in_buf[733]*(4)+in_buf[734]*(28)+in_buf[735]*(32)+in_buf[736]*(13)+in_buf[737]*(24)+in_buf[738]*(32)+in_buf[739]*(5)+in_buf[740]*(-1)+in_buf[741]*(7)+in_buf[742]*(36)+in_buf[743]*(32)+in_buf[744]*(29)+in_buf[745]*(23)+in_buf[746]*(2)+in_buf[747]*(0)+in_buf[748]*(23)+in_buf[749]*(10)+in_buf[750]*(9)+in_buf[751]*(-11)+in_buf[752]*(6)+in_buf[753]*(8)+in_buf[754]*(2)+in_buf[755]*(0)+in_buf[756]*(-1)+in_buf[757]*(-3)+in_buf[758]*(1)+in_buf[759]*(0)+in_buf[760]*(-19)+in_buf[761]*(-15)+in_buf[762]*(15)+in_buf[763]*(12)+in_buf[764]*(19)+in_buf[765]*(11)+in_buf[766]*(48)+in_buf[767]*(31)+in_buf[768]*(26)+in_buf[769]*(29)+in_buf[770]*(70)+in_buf[771]*(52)+in_buf[772]*(46)+in_buf[773]*(34)+in_buf[774]*(12)+in_buf[775]*(19)+in_buf[776]*(27)+in_buf[777]*(29)+in_buf[778]*(25)+in_buf[779]*(20)+in_buf[780]*(4)+in_buf[781]*(3)+in_buf[782]*(0)+in_buf[783]*(-1);
assign in_buf_weight023=in_buf[0]*(0)+in_buf[1]*(1)+in_buf[2]*(0)+in_buf[3]*(3)+in_buf[4]*(1)+in_buf[5]*(2)+in_buf[6]*(-1)+in_buf[7]*(-2)+in_buf[8]*(1)+in_buf[9]*(-3)+in_buf[10]*(0)+in_buf[11]*(1)+in_buf[12]*(-10)+in_buf[13]*(-10)+in_buf[14]*(7)+in_buf[15]*(6)+in_buf[16]*(0)+in_buf[17]*(-3)+in_buf[18]*(3)+in_buf[19]*(0)+in_buf[20]*(-3)+in_buf[21]*(3)+in_buf[22]*(-2)+in_buf[23]*(0)+in_buf[24]*(3)+in_buf[25]*(0)+in_buf[26]*(0)+in_buf[27]*(4)+in_buf[28]*(4)+in_buf[29]*(-4)+in_buf[30]*(3)+in_buf[31]*(-1)+in_buf[32]*(-9)+in_buf[33]*(-11)+in_buf[34]*(-2)+in_buf[35]*(-5)+in_buf[36]*(-11)+in_buf[37]*(-5)+in_buf[38]*(-10)+in_buf[39]*(-11)+in_buf[40]*(-13)+in_buf[41]*(-25)+in_buf[42]*(21)+in_buf[43]*(20)+in_buf[44]*(10)+in_buf[45]*(-3)+in_buf[46]*(-10)+in_buf[47]*(-11)+in_buf[48]*(-29)+in_buf[49]*(-19)+in_buf[50]*(-2)+in_buf[51]*(-1)+in_buf[52]*(1)+in_buf[53]*(-3)+in_buf[54]*(1)+in_buf[55]*(0)+in_buf[56]*(-2)+in_buf[57]*(0)+in_buf[58]*(-15)+in_buf[59]*(1)+in_buf[60]*(-10)+in_buf[61]*(-6)+in_buf[62]*(-15)+in_buf[63]*(-19)+in_buf[64]*(-19)+in_buf[65]*(13)+in_buf[66]*(18)+in_buf[67]*(2)+in_buf[68]*(3)+in_buf[69]*(25)+in_buf[70]*(7)+in_buf[71]*(17)+in_buf[72]*(23)+in_buf[73]*(12)+in_buf[74]*(4)+in_buf[75]*(8)+in_buf[76]*(7)+in_buf[77]*(-9)+in_buf[78]*(-14)+in_buf[79]*(6)+in_buf[80]*(9)+in_buf[81]*(7)+in_buf[82]*(-2)+in_buf[83]*(-3)+in_buf[84]*(0)+in_buf[85]*(2)+in_buf[86]*(14)+in_buf[87]*(20)+in_buf[88]*(3)+in_buf[89]*(-5)+in_buf[90]*(-5)+in_buf[91]*(-4)+in_buf[92]*(18)+in_buf[93]*(4)+in_buf[94]*(28)+in_buf[95]*(4)+in_buf[96]*(7)+in_buf[97]*(2)+in_buf[98]*(-14)+in_buf[99]*(16)+in_buf[100]*(40)+in_buf[101]*(22)+in_buf[102]*(28)+in_buf[103]*(21)+in_buf[104]*(13)+in_buf[105]*(-4)+in_buf[106]*(-7)+in_buf[107]*(5)+in_buf[108]*(8)+in_buf[109]*(7)+in_buf[110]*(-21)+in_buf[111]*(0)+in_buf[112]*(3)+in_buf[113]*(2)+in_buf[114]*(13)+in_buf[115]*(-1)+in_buf[116]*(3)+in_buf[117]*(20)+in_buf[118]*(12)+in_buf[119]*(20)+in_buf[120]*(34)+in_buf[121]*(27)+in_buf[122]*(36)+in_buf[123]*(44)+in_buf[124]*(38)+in_buf[125]*(24)+in_buf[126]*(14)+in_buf[127]*(33)+in_buf[128]*(46)+in_buf[129]*(26)+in_buf[130]*(25)+in_buf[131]*(29)+in_buf[132]*(16)+in_buf[133]*(3)+in_buf[134]*(9)+in_buf[135]*(-11)+in_buf[136]*(3)+in_buf[137]*(-5)+in_buf[138]*(-7)+in_buf[139]*(-15)+in_buf[140]*(1)+in_buf[141]*(4)+in_buf[142]*(14)+in_buf[143]*(38)+in_buf[144]*(53)+in_buf[145]*(23)+in_buf[146]*(21)+in_buf[147]*(18)+in_buf[148]*(-2)+in_buf[149]*(14)+in_buf[150]*(18)+in_buf[151]*(14)+in_buf[152]*(11)+in_buf[153]*(-2)+in_buf[154]*(-4)+in_buf[155]*(12)+in_buf[156]*(15)+in_buf[157]*(3)+in_buf[158]*(6)+in_buf[159]*(19)+in_buf[160]*(25)+in_buf[161]*(6)+in_buf[162]*(13)+in_buf[163]*(-7)+in_buf[164]*(-9)+in_buf[165]*(-3)+in_buf[166]*(-14)+in_buf[167]*(-18)+in_buf[168]*(1)+in_buf[169]*(3)+in_buf[170]*(-25)+in_buf[171]*(7)+in_buf[172]*(3)+in_buf[173]*(-8)+in_buf[174]*(20)+in_buf[175]*(7)+in_buf[176]*(11)+in_buf[177]*(14)+in_buf[178]*(20)+in_buf[179]*(15)+in_buf[180]*(6)+in_buf[181]*(2)+in_buf[182]*(7)+in_buf[183]*(0)+in_buf[184]*(2)+in_buf[185]*(-7)+in_buf[186]*(-1)+in_buf[187]*(-12)+in_buf[188]*(2)+in_buf[189]*(-11)+in_buf[190]*(-14)+in_buf[191]*(-9)+in_buf[192]*(-28)+in_buf[193]*(-9)+in_buf[194]*(6)+in_buf[195]*(-19)+in_buf[196]*(-11)+in_buf[197]*(-1)+in_buf[198]*(-31)+in_buf[199]*(-10)+in_buf[200]*(16)+in_buf[201]*(-11)+in_buf[202]*(16)+in_buf[203]*(12)+in_buf[204]*(13)+in_buf[205]*(-3)+in_buf[206]*(10)+in_buf[207]*(-5)+in_buf[208]*(7)+in_buf[209]*(15)+in_buf[210]*(6)+in_buf[211]*(-2)+in_buf[212]*(1)+in_buf[213]*(-13)+in_buf[214]*(-9)+in_buf[215]*(-11)+in_buf[216]*(-11)+in_buf[217]*(-13)+in_buf[218]*(0)+in_buf[219]*(-5)+in_buf[220]*(-18)+in_buf[221]*(9)+in_buf[222]*(0)+in_buf[223]*(-25)+in_buf[224]*(1)+in_buf[225]*(-29)+in_buf[226]*(-27)+in_buf[227]*(24)+in_buf[228]*(9)+in_buf[229]*(-5)+in_buf[230]*(4)+in_buf[231]*(6)+in_buf[232]*(-9)+in_buf[233]*(-22)+in_buf[234]*(-9)+in_buf[235]*(-4)+in_buf[236]*(5)+in_buf[237]*(13)+in_buf[238]*(-1)+in_buf[239]*(2)+in_buf[240]*(-1)+in_buf[241]*(-1)+in_buf[242]*(4)+in_buf[243]*(7)+in_buf[244]*(-6)+in_buf[245]*(-12)+in_buf[246]*(8)+in_buf[247]*(12)+in_buf[248]*(-19)+in_buf[249]*(17)+in_buf[250]*(39)+in_buf[251]*(20)+in_buf[252]*(-13)+in_buf[253]*(-25)+in_buf[254]*(4)+in_buf[255]*(32)+in_buf[256]*(-3)+in_buf[257]*(-16)+in_buf[258]*(-14)+in_buf[259]*(-6)+in_buf[260]*(0)+in_buf[261]*(-10)+in_buf[262]*(14)+in_buf[263]*(13)+in_buf[264]*(7)+in_buf[265]*(-2)+in_buf[266]*(-8)+in_buf[267]*(11)+in_buf[268]*(3)+in_buf[269]*(3)+in_buf[270]*(6)+in_buf[271]*(11)+in_buf[272]*(-6)+in_buf[273]*(-6)+in_buf[274]*(20)+in_buf[275]*(14)+in_buf[276]*(-18)+in_buf[277]*(23)+in_buf[278]*(44)+in_buf[279]*(20)+in_buf[280]*(-10)+in_buf[281]*(-11)+in_buf[282]*(-11)+in_buf[283]*(21)+in_buf[284]*(-11)+in_buf[285]*(-34)+in_buf[286]*(-16)+in_buf[287]*(-7)+in_buf[288]*(-11)+in_buf[289]*(-21)+in_buf[290]*(13)+in_buf[291]*(9)+in_buf[292]*(14)+in_buf[293]*(-4)+in_buf[294]*(2)+in_buf[295]*(0)+in_buf[296]*(14)+in_buf[297]*(16)+in_buf[298]*(16)+in_buf[299]*(5)+in_buf[300]*(-12)+in_buf[301]*(-14)+in_buf[302]*(5)+in_buf[303]*(5)+in_buf[304]*(-30)+in_buf[305]*(1)+in_buf[306]*(29)+in_buf[307]*(32)+in_buf[308]*(-14)+in_buf[309]*(-14)+in_buf[310]*(-22)+in_buf[311]*(-5)+in_buf[312]*(-17)+in_buf[313]*(-38)+in_buf[314]*(-34)+in_buf[315]*(-15)+in_buf[316]*(-42)+in_buf[317]*(-44)+in_buf[318]*(-8)+in_buf[319]*(1)+in_buf[320]*(0)+in_buf[321]*(-4)+in_buf[322]*(4)+in_buf[323]*(16)+in_buf[324]*(22)+in_buf[325]*(33)+in_buf[326]*(21)+in_buf[327]*(3)+in_buf[328]*(-16)+in_buf[329]*(-30)+in_buf[330]*(-25)+in_buf[331]*(-22)+in_buf[332]*(-25)+in_buf[333]*(9)+in_buf[334]*(33)+in_buf[335]*(27)+in_buf[336]*(-23)+in_buf[337]*(-14)+in_buf[338]*(-7)+in_buf[339]*(-2)+in_buf[340]*(-28)+in_buf[341]*(-43)+in_buf[342]*(-35)+in_buf[343]*(-30)+in_buf[344]*(-36)+in_buf[345]*(-18)+in_buf[346]*(-10)+in_buf[347]*(-9)+in_buf[348]*(-3)+in_buf[349]*(3)+in_buf[350]*(24)+in_buf[351]*(30)+in_buf[352]*(32)+in_buf[353]*(31)+in_buf[354]*(9)+in_buf[355]*(-6)+in_buf[356]*(-29)+in_buf[357]*(-33)+in_buf[358]*(-39)+in_buf[359]*(-22)+in_buf[360]*(-31)+in_buf[361]*(-12)+in_buf[362]*(16)+in_buf[363]*(19)+in_buf[364]*(20)+in_buf[365]*(-8)+in_buf[366]*(-35)+in_buf[367]*(-18)+in_buf[368]*(-35)+in_buf[369]*(-49)+in_buf[370]*(-36)+in_buf[371]*(-12)+in_buf[372]*(-15)+in_buf[373]*(-11)+in_buf[374]*(-12)+in_buf[375]*(6)+in_buf[376]*(11)+in_buf[377]*(22)+in_buf[378]*(37)+in_buf[379]*(29)+in_buf[380]*(30)+in_buf[381]*(21)+in_buf[382]*(-3)+in_buf[383]*(-32)+in_buf[384]*(-28)+in_buf[385]*(-24)+in_buf[386]*(-9)+in_buf[387]*(-12)+in_buf[388]*(-19)+in_buf[389]*(-26)+in_buf[390]*(23)+in_buf[391]*(2)+in_buf[392]*(-20)+in_buf[393]*(0)+in_buf[394]*(-9)+in_buf[395]*(-8)+in_buf[396]*(-15)+in_buf[397]*(-39)+in_buf[398]*(-16)+in_buf[399]*(-5)+in_buf[400]*(-11)+in_buf[401]*(-7)+in_buf[402]*(-14)+in_buf[403]*(-15)+in_buf[404]*(-5)+in_buf[405]*(16)+in_buf[406]*(32)+in_buf[407]*(10)+in_buf[408]*(9)+in_buf[409]*(-4)+in_buf[410]*(-15)+in_buf[411]*(-36)+in_buf[412]*(-31)+in_buf[413]*(-11)+in_buf[414]*(0)+in_buf[415]*(-10)+in_buf[416]*(9)+in_buf[417]*(-11)+in_buf[418]*(38)+in_buf[419]*(3)+in_buf[420]*(-14)+in_buf[421]*(7)+in_buf[422]*(14)+in_buf[423]*(5)+in_buf[424]*(12)+in_buf[425]*(-15)+in_buf[426]*(-8)+in_buf[427]*(-14)+in_buf[428]*(-7)+in_buf[429]*(0)+in_buf[430]*(-16)+in_buf[431]*(-5)+in_buf[432]*(-11)+in_buf[433]*(19)+in_buf[434]*(12)+in_buf[435]*(-5)+in_buf[436]*(-8)+in_buf[437]*(-27)+in_buf[438]*(-35)+in_buf[439]*(-24)+in_buf[440]*(-20)+in_buf[441]*(-17)+in_buf[442]*(-12)+in_buf[443]*(-10)+in_buf[444]*(15)+in_buf[445]*(23)+in_buf[446]*(25)+in_buf[447]*(21)+in_buf[448]*(1)+in_buf[449]*(28)+in_buf[450]*(15)+in_buf[451]*(23)+in_buf[452]*(13)+in_buf[453]*(-3)+in_buf[454]*(7)+in_buf[455]*(-14)+in_buf[456]*(-19)+in_buf[457]*(-4)+in_buf[458]*(-7)+in_buf[459]*(-25)+in_buf[460]*(-12)+in_buf[461]*(3)+in_buf[462]*(11)+in_buf[463]*(-11)+in_buf[464]*(-15)+in_buf[465]*(-35)+in_buf[466]*(-15)+in_buf[467]*(-9)+in_buf[468]*(-8)+in_buf[469]*(5)+in_buf[470]*(6)+in_buf[471]*(1)+in_buf[472]*(18)+in_buf[473]*(53)+in_buf[474]*(35)+in_buf[475]*(23)+in_buf[476]*(-3)+in_buf[477]*(14)+in_buf[478]*(11)+in_buf[479]*(41)+in_buf[480]*(13)+in_buf[481]*(14)+in_buf[482]*(10)+in_buf[483]*(-1)+in_buf[484]*(0)+in_buf[485]*(-1)+in_buf[486]*(-8)+in_buf[487]*(-29)+in_buf[488]*(-16)+in_buf[489]*(10)+in_buf[490]*(17)+in_buf[491]*(1)+in_buf[492]*(-7)+in_buf[493]*(-11)+in_buf[494]*(-9)+in_buf[495]*(4)+in_buf[496]*(1)+in_buf[497]*(7)+in_buf[498]*(-1)+in_buf[499]*(4)+in_buf[500]*(22)+in_buf[501]*(39)+in_buf[502]*(29)+in_buf[503]*(38)+in_buf[504]*(-31)+in_buf[505]*(17)+in_buf[506]*(26)+in_buf[507]*(43)+in_buf[508]*(15)+in_buf[509]*(31)+in_buf[510]*(21)+in_buf[511]*(-2)+in_buf[512]*(8)+in_buf[513]*(15)+in_buf[514]*(0)+in_buf[515]*(-12)+in_buf[516]*(-29)+in_buf[517]*(1)+in_buf[518]*(7)+in_buf[519]*(-3)+in_buf[520]*(15)+in_buf[521]*(16)+in_buf[522]*(1)+in_buf[523]*(13)+in_buf[524]*(9)+in_buf[525]*(0)+in_buf[526]*(1)+in_buf[527]*(14)+in_buf[528]*(32)+in_buf[529]*(41)+in_buf[530]*(11)+in_buf[531]*(16)+in_buf[532]*(23)+in_buf[533]*(-10)+in_buf[534]*(-10)+in_buf[535]*(4)+in_buf[536]*(25)+in_buf[537]*(31)+in_buf[538]*(20)+in_buf[539]*(12)+in_buf[540]*(16)+in_buf[541]*(24)+in_buf[542]*(12)+in_buf[543]*(-9)+in_buf[544]*(-18)+in_buf[545]*(6)+in_buf[546]*(-8)+in_buf[547]*(8)+in_buf[548]*(28)+in_buf[549]*(17)+in_buf[550]*(9)+in_buf[551]*(12)+in_buf[552]*(0)+in_buf[553]*(2)+in_buf[554]*(-7)+in_buf[555]*(6)+in_buf[556]*(27)+in_buf[557]*(55)+in_buf[558]*(40)+in_buf[559]*(-2)+in_buf[560]*(-1)+in_buf[561]*(-2)+in_buf[562]*(-4)+in_buf[563]*(9)+in_buf[564]*(28)+in_buf[565]*(27)+in_buf[566]*(29)+in_buf[567]*(12)+in_buf[568]*(12)+in_buf[569]*(13)+in_buf[570]*(11)+in_buf[571]*(-1)+in_buf[572]*(-11)+in_buf[573]*(-8)+in_buf[574]*(-7)+in_buf[575]*(4)+in_buf[576]*(20)+in_buf[577]*(19)+in_buf[578]*(14)+in_buf[579]*(21)+in_buf[580]*(13)+in_buf[581]*(6)+in_buf[582]*(-7)+in_buf[583]*(7)+in_buf[584]*(4)+in_buf[585]*(7)+in_buf[586]*(24)+in_buf[587]*(17)+in_buf[588]*(19)+in_buf[589]*(1)+in_buf[590]*(33)+in_buf[591]*(15)+in_buf[592]*(12)+in_buf[593]*(3)+in_buf[594]*(9)+in_buf[595]*(1)+in_buf[596]*(6)+in_buf[597]*(6)+in_buf[598]*(9)+in_buf[599]*(-2)+in_buf[600]*(-6)+in_buf[601]*(-10)+in_buf[602]*(-13)+in_buf[603]*(-5)+in_buf[604]*(7)+in_buf[605]*(-3)+in_buf[606]*(22)+in_buf[607]*(22)+in_buf[608]*(16)+in_buf[609]*(6)+in_buf[610]*(3)+in_buf[611]*(13)+in_buf[612]*(7)+in_buf[613]*(18)+in_buf[614]*(-25)+in_buf[615]*(-4)+in_buf[616]*(14)+in_buf[617]*(11)+in_buf[618]*(17)+in_buf[619]*(27)+in_buf[620]*(26)+in_buf[621]*(21)+in_buf[622]*(-4)+in_buf[623]*(0)+in_buf[624]*(1)+in_buf[625]*(0)+in_buf[626]*(-3)+in_buf[627]*(-2)+in_buf[628]*(-11)+in_buf[629]*(-6)+in_buf[630]*(1)+in_buf[631]*(-6)+in_buf[632]*(-1)+in_buf[633]*(11)+in_buf[634]*(23)+in_buf[635]*(12)+in_buf[636]*(39)+in_buf[637]*(7)+in_buf[638]*(-4)+in_buf[639]*(-3)+in_buf[640]*(27)+in_buf[641]*(30)+in_buf[642]*(-2)+in_buf[643]*(1)+in_buf[644]*(2)+in_buf[645]*(-3)+in_buf[646]*(13)+in_buf[647]*(13)+in_buf[648]*(12)+in_buf[649]*(2)+in_buf[650]*(-12)+in_buf[651]*(-10)+in_buf[652]*(11)+in_buf[653]*(8)+in_buf[654]*(0)+in_buf[655]*(0)+in_buf[656]*(-1)+in_buf[657]*(-5)+in_buf[658]*(-4)+in_buf[659]*(9)+in_buf[660]*(10)+in_buf[661]*(18)+in_buf[662]*(21)+in_buf[663]*(23)+in_buf[664]*(35)+in_buf[665]*(17)+in_buf[666]*(27)+in_buf[667]*(30)+in_buf[668]*(13)+in_buf[669]*(24)+in_buf[670]*(29)+in_buf[671]*(1)+in_buf[672]*(0)+in_buf[673]*(3)+in_buf[674]*(5)+in_buf[675]*(-1)+in_buf[676]*(5)+in_buf[677]*(-9)+in_buf[678]*(-10)+in_buf[679]*(0)+in_buf[680]*(0)+in_buf[681]*(-2)+in_buf[682]*(10)+in_buf[683]*(2)+in_buf[684]*(-14)+in_buf[685]*(-23)+in_buf[686]*(-21)+in_buf[687]*(-10)+in_buf[688]*(-1)+in_buf[689]*(12)+in_buf[690]*(14)+in_buf[691]*(6)+in_buf[692]*(0)+in_buf[693]*(2)+in_buf[694]*(-4)+in_buf[695]*(12)+in_buf[696]*(25)+in_buf[697]*(27)+in_buf[698]*(15)+in_buf[699]*(0)+in_buf[700]*(-2)+in_buf[701]*(-1)+in_buf[702]*(5)+in_buf[703]*(-21)+in_buf[704]*(-26)+in_buf[705]*(-22)+in_buf[706]*(-2)+in_buf[707]*(-8)+in_buf[708]*(20)+in_buf[709]*(22)+in_buf[710]*(-5)+in_buf[711]*(-22)+in_buf[712]*(13)+in_buf[713]*(15)+in_buf[714]*(28)+in_buf[715]*(17)+in_buf[716]*(39)+in_buf[717]*(47)+in_buf[718]*(14)+in_buf[719]*(-8)+in_buf[720]*(-14)+in_buf[721]*(-13)+in_buf[722]*(-21)+in_buf[723]*(-29)+in_buf[724]*(-4)+in_buf[725]*(14)+in_buf[726]*(5)+in_buf[727]*(2)+in_buf[728]*(3)+in_buf[729]*(-2)+in_buf[730]*(0)+in_buf[731]*(7)+in_buf[732]*(14)+in_buf[733]*(-25)+in_buf[734]*(-43)+in_buf[735]*(-28)+in_buf[736]*(-5)+in_buf[737]*(16)+in_buf[738]*(14)+in_buf[739]*(-6)+in_buf[740]*(-16)+in_buf[741]*(-7)+in_buf[742]*(23)+in_buf[743]*(34)+in_buf[744]*(44)+in_buf[745]*(60)+in_buf[746]*(27)+in_buf[747]*(-6)+in_buf[748]*(10)+in_buf[749]*(17)+in_buf[750]*(14)+in_buf[751]*(-1)+in_buf[752]*(7)+in_buf[753]*(-6)+in_buf[754]*(1)+in_buf[755]*(4)+in_buf[756]*(0)+in_buf[757]*(3)+in_buf[758]*(-1)+in_buf[759]*(3)+in_buf[760]*(-12)+in_buf[761]*(-6)+in_buf[762]*(-12)+in_buf[763]*(-18)+in_buf[764]*(-1)+in_buf[765]*(7)+in_buf[766]*(-7)+in_buf[767]*(4)+in_buf[768]*(5)+in_buf[769]*(24)+in_buf[770]*(54)+in_buf[771]*(42)+in_buf[772]*(1)+in_buf[773]*(-5)+in_buf[774]*(28)+in_buf[775]*(4)+in_buf[776]*(-8)+in_buf[777]*(7)+in_buf[778]*(-1)+in_buf[779]*(-2)+in_buf[780]*(0)+in_buf[781]*(4)+in_buf[782]*(2)+in_buf[783]*(-1);
assign in_buf_weight024=in_buf[0]*(-2)+in_buf[1]*(-1)+in_buf[2]*(1)+in_buf[3]*(-2)+in_buf[4]*(2)+in_buf[5]*(1)+in_buf[6]*(0)+in_buf[7]*(2)+in_buf[8]*(1)+in_buf[9]*(-2)+in_buf[10]*(-3)+in_buf[11]*(1)+in_buf[12]*(7)+in_buf[13]*(6)+in_buf[14]*(-19)+in_buf[15]*(-15)+in_buf[16]*(-1)+in_buf[17]*(-1)+in_buf[18]*(0)+in_buf[19]*(4)+in_buf[20]*(3)+in_buf[21]*(3)+in_buf[22]*(4)+in_buf[23]*(0)+in_buf[24]*(0)+in_buf[25]*(2)+in_buf[26]*(-3)+in_buf[27]*(3)+in_buf[28]*(-1)+in_buf[29]*(-3)+in_buf[30]*(0)+in_buf[31]*(2)+in_buf[32]*(7)+in_buf[33]*(-4)+in_buf[34]*(-2)+in_buf[35]*(-4)+in_buf[36]*(17)+in_buf[37]*(15)+in_buf[38]*(17)+in_buf[39]*(1)+in_buf[40]*(5)+in_buf[41]*(28)+in_buf[42]*(1)+in_buf[43]*(-22)+in_buf[44]*(-10)+in_buf[45]*(12)+in_buf[46]*(25)+in_buf[47]*(18)+in_buf[48]*(29)+in_buf[49]*(29)+in_buf[50]*(18)+in_buf[51]*(15)+in_buf[52]*(0)+in_buf[53]*(3)+in_buf[54]*(4)+in_buf[55]*(-1)+in_buf[56]*(1)+in_buf[57]*(-2)+in_buf[58]*(8)+in_buf[59]*(-30)+in_buf[60]*(-16)+in_buf[61]*(9)+in_buf[62]*(10)+in_buf[63]*(20)+in_buf[64]*(18)+in_buf[65]*(-5)+in_buf[66]*(-5)+in_buf[67]*(22)+in_buf[68]*(0)+in_buf[69]*(-28)+in_buf[70]*(0)+in_buf[71]*(-9)+in_buf[72]*(-19)+in_buf[73]*(-7)+in_buf[74]*(-3)+in_buf[75]*(-4)+in_buf[76]*(0)+in_buf[77]*(8)+in_buf[78]*(26)+in_buf[79]*(1)+in_buf[80]*(-5)+in_buf[81]*(-11)+in_buf[82]*(4)+in_buf[83]*(-1)+in_buf[84]*(-1)+in_buf[85]*(3)+in_buf[86]*(-14)+in_buf[87]*(-31)+in_buf[88]*(-8)+in_buf[89]*(6)+in_buf[90]*(0)+in_buf[91]*(19)+in_buf[92]*(-10)+in_buf[93]*(-6)+in_buf[94]*(-5)+in_buf[95]*(10)+in_buf[96]*(0)+in_buf[97]*(5)+in_buf[98]*(2)+in_buf[99]*(0)+in_buf[100]*(-13)+in_buf[101]*(2)+in_buf[102]*(12)+in_buf[103]*(-3)+in_buf[104]*(4)+in_buf[105]*(33)+in_buf[106]*(33)+in_buf[107]*(33)+in_buf[108]*(11)+in_buf[109]*(-5)+in_buf[110]*(2)+in_buf[111]*(4)+in_buf[112]*(-3)+in_buf[113]*(-5)+in_buf[114]*(-16)+in_buf[115]*(-10)+in_buf[116]*(14)+in_buf[117]*(-16)+in_buf[118]*(3)+in_buf[119]*(19)+in_buf[120]*(-19)+in_buf[121]*(-12)+in_buf[122]*(1)+in_buf[123]*(-7)+in_buf[124]*(0)+in_buf[125]*(-7)+in_buf[126]*(-2)+in_buf[127]*(-6)+in_buf[128]*(-1)+in_buf[129]*(12)+in_buf[130]*(8)+in_buf[131]*(5)+in_buf[132]*(13)+in_buf[133]*(9)+in_buf[134]*(7)+in_buf[135]*(24)+in_buf[136]*(11)+in_buf[137]*(4)+in_buf[138]*(-18)+in_buf[139]*(4)+in_buf[140]*(4)+in_buf[141]*(3)+in_buf[142]*(-11)+in_buf[143]*(-16)+in_buf[144]*(-14)+in_buf[145]*(-37)+in_buf[146]*(-23)+in_buf[147]*(-9)+in_buf[148]*(-13)+in_buf[149]*(4)+in_buf[150]*(10)+in_buf[151]*(18)+in_buf[152]*(16)+in_buf[153]*(12)+in_buf[154]*(13)+in_buf[155]*(20)+in_buf[156]*(23)+in_buf[157]*(20)+in_buf[158]*(5)+in_buf[159]*(-2)+in_buf[160]*(8)+in_buf[161]*(3)+in_buf[162]*(-30)+in_buf[163]*(-21)+in_buf[164]*(1)+in_buf[165]*(-3)+in_buf[166]*(0)+in_buf[167]*(3)+in_buf[168]*(0)+in_buf[169]*(-11)+in_buf[170]*(-7)+in_buf[171]*(-21)+in_buf[172]*(8)+in_buf[173]*(-17)+in_buf[174]*(-19)+in_buf[175]*(0)+in_buf[176]*(-1)+in_buf[177]*(-1)+in_buf[178]*(0)+in_buf[179]*(0)+in_buf[180]*(3)+in_buf[181]*(7)+in_buf[182]*(14)+in_buf[183]*(13)+in_buf[184]*(13)+in_buf[185]*(0)+in_buf[186]*(-13)+in_buf[187]*(-4)+in_buf[188]*(7)+in_buf[189]*(-9)+in_buf[190]*(-20)+in_buf[191]*(-2)+in_buf[192]*(12)+in_buf[193]*(5)+in_buf[194]*(-16)+in_buf[195]*(3)+in_buf[196]*(1)+in_buf[197]*(-29)+in_buf[198]*(-1)+in_buf[199]*(-30)+in_buf[200]*(-20)+in_buf[201]*(0)+in_buf[202]*(-1)+in_buf[203]*(-12)+in_buf[204]*(-9)+in_buf[205]*(0)+in_buf[206]*(-6)+in_buf[207]*(-5)+in_buf[208]*(-11)+in_buf[209]*(5)+in_buf[210]*(1)+in_buf[211]*(6)+in_buf[212]*(-6)+in_buf[213]*(-3)+in_buf[214]*(-21)+in_buf[215]*(-11)+in_buf[216]*(-7)+in_buf[217]*(0)+in_buf[218]*(-10)+in_buf[219]*(-11)+in_buf[220]*(24)+in_buf[221]*(22)+in_buf[222]*(3)+in_buf[223]*(7)+in_buf[224]*(-19)+in_buf[225]*(-11)+in_buf[226]*(5)+in_buf[227]*(-10)+in_buf[228]*(5)+in_buf[229]*(10)+in_buf[230]*(9)+in_buf[231]*(-16)+in_buf[232]*(-10)+in_buf[233]*(-7)+in_buf[234]*(-14)+in_buf[235]*(-5)+in_buf[236]*(-17)+in_buf[237]*(-16)+in_buf[238]*(0)+in_buf[239]*(0)+in_buf[240]*(-4)+in_buf[241]*(-15)+in_buf[242]*(-13)+in_buf[243]*(-5)+in_buf[244]*(-5)+in_buf[245]*(15)+in_buf[246]*(-26)+in_buf[247]*(-35)+in_buf[248]*(42)+in_buf[249]*(39)+in_buf[250]*(4)+in_buf[251]*(-20)+in_buf[252]*(0)+in_buf[253]*(-9)+in_buf[254]*(-7)+in_buf[255]*(-13)+in_buf[256]*(-7)+in_buf[257]*(0)+in_buf[258]*(18)+in_buf[259]*(-10)+in_buf[260]*(-19)+in_buf[261]*(-4)+in_buf[262]*(-3)+in_buf[263]*(0)+in_buf[264]*(-21)+in_buf[265]*(-12)+in_buf[266]*(-17)+in_buf[267]*(-10)+in_buf[268]*(-12)+in_buf[269]*(-10)+in_buf[270]*(-11)+in_buf[271]*(-5)+in_buf[272]*(8)+in_buf[273]*(6)+in_buf[274]*(-32)+in_buf[275]*(-23)+in_buf[276]*(24)+in_buf[277]*(-11)+in_buf[278]*(-7)+in_buf[279]*(-18)+in_buf[280]*(-1)+in_buf[281]*(-7)+in_buf[282]*(-25)+in_buf[283]*(1)+in_buf[284]*(-25)+in_buf[285]*(6)+in_buf[286]*(9)+in_buf[287]*(-2)+in_buf[288]*(-14)+in_buf[289]*(-3)+in_buf[290]*(0)+in_buf[291]*(-11)+in_buf[292]*(-26)+in_buf[293]*(-35)+in_buf[294]*(-24)+in_buf[295]*(-21)+in_buf[296]*(-26)+in_buf[297]*(-17)+in_buf[298]*(-7)+in_buf[299]*(-5)+in_buf[300]*(-6)+in_buf[301]*(-6)+in_buf[302]*(-22)+in_buf[303]*(-4)+in_buf[304]*(7)+in_buf[305]*(-7)+in_buf[306]*(-16)+in_buf[307]*(-15)+in_buf[308]*(-1)+in_buf[309]*(-33)+in_buf[310]*(-30)+in_buf[311]*(-15)+in_buf[312]*(-26)+in_buf[313]*(6)+in_buf[314]*(23)+in_buf[315]*(0)+in_buf[316]*(9)+in_buf[317]*(19)+in_buf[318]*(18)+in_buf[319]*(-9)+in_buf[320]*(-31)+in_buf[321]*(-26)+in_buf[322]*(-9)+in_buf[323]*(-7)+in_buf[324]*(-4)+in_buf[325]*(4)+in_buf[326]*(-3)+in_buf[327]*(1)+in_buf[328]*(-11)+in_buf[329]*(-4)+in_buf[330]*(2)+in_buf[331]*(-8)+in_buf[332]*(-14)+in_buf[333]*(-27)+in_buf[334]*(-8)+in_buf[335]*(-31)+in_buf[336]*(-1)+in_buf[337]*(-1)+in_buf[338]*(-4)+in_buf[339]*(-9)+in_buf[340]*(1)+in_buf[341]*(19)+in_buf[342]*(33)+in_buf[343]*(14)+in_buf[344]*(11)+in_buf[345]*(24)+in_buf[346]*(18)+in_buf[347]*(-1)+in_buf[348]*(-28)+in_buf[349]*(-25)+in_buf[350]*(-10)+in_buf[351]*(-4)+in_buf[352]*(-13)+in_buf[353]*(15)+in_buf[354]*(4)+in_buf[355]*(13)+in_buf[356]*(6)+in_buf[357]*(12)+in_buf[358]*(24)+in_buf[359]*(27)+in_buf[360]*(-7)+in_buf[361]*(-37)+in_buf[362]*(-21)+in_buf[363]*(-37)+in_buf[364]*(-3)+in_buf[365]*(0)+in_buf[366]*(-13)+in_buf[367]*(0)+in_buf[368]*(32)+in_buf[369]*(34)+in_buf[370]*(29)+in_buf[371]*(31)+in_buf[372]*(23)+in_buf[373]*(28)+in_buf[374]*(41)+in_buf[375]*(-5)+in_buf[376]*(-18)+in_buf[377]*(-9)+in_buf[378]*(0)+in_buf[379]*(2)+in_buf[380]*(-5)+in_buf[381]*(0)+in_buf[382]*(21)+in_buf[383]*(30)+in_buf[384]*(14)+in_buf[385]*(18)+in_buf[386]*(26)+in_buf[387]*(37)+in_buf[388]*(0)+in_buf[389]*(-27)+in_buf[390]*(-26)+in_buf[391]*(-14)+in_buf[392]*(0)+in_buf[393]*(-6)+in_buf[394]*(-21)+in_buf[395]*(13)+in_buf[396]*(34)+in_buf[397]*(31)+in_buf[398]*(25)+in_buf[399]*(25)+in_buf[400]*(17)+in_buf[401]*(29)+in_buf[402]*(19)+in_buf[403]*(8)+in_buf[404]*(9)+in_buf[405]*(4)+in_buf[406]*(-1)+in_buf[407]*(-1)+in_buf[408]*(2)+in_buf[409]*(6)+in_buf[410]*(14)+in_buf[411]*(20)+in_buf[412]*(31)+in_buf[413]*(21)+in_buf[414]*(11)+in_buf[415]*(6)+in_buf[416]*(-14)+in_buf[417]*(6)+in_buf[418]*(-20)+in_buf[419]*(-9)+in_buf[420]*(-3)+in_buf[421]*(-11)+in_buf[422]*(2)+in_buf[423]*(28)+in_buf[424]*(21)+in_buf[425]*(9)+in_buf[426]*(9)+in_buf[427]*(21)+in_buf[428]*(13)+in_buf[429]*(11)+in_buf[430]*(19)+in_buf[431]*(11)+in_buf[432]*(22)+in_buf[433]*(14)+in_buf[434]*(-6)+in_buf[435]*(-7)+in_buf[436]*(0)+in_buf[437]*(11)+in_buf[438]*(11)+in_buf[439]*(28)+in_buf[440]*(24)+in_buf[441]*(13)+in_buf[442]*(12)+in_buf[443]*(-6)+in_buf[444]*(-38)+in_buf[445]*(22)+in_buf[446]*(5)+in_buf[447]*(-11)+in_buf[448]*(-6)+in_buf[449]*(-10)+in_buf[450]*(3)+in_buf[451]*(7)+in_buf[452]*(-8)+in_buf[453]*(8)+in_buf[454]*(14)+in_buf[455]*(15)+in_buf[456]*(24)+in_buf[457]*(1)+in_buf[458]*(11)+in_buf[459]*(27)+in_buf[460]*(30)+in_buf[461]*(0)+in_buf[462]*(-3)+in_buf[463]*(0)+in_buf[464]*(2)+in_buf[465]*(16)+in_buf[466]*(25)+in_buf[467]*(15)+in_buf[468]*(24)+in_buf[469]*(1)+in_buf[470]*(13)+in_buf[471]*(1)+in_buf[472]*(-22)+in_buf[473]*(34)+in_buf[474]*(-10)+in_buf[475]*(-20)+in_buf[476]*(0)+in_buf[477]*(-3)+in_buf[478]*(6)+in_buf[479]*(-4)+in_buf[480]*(-18)+in_buf[481]*(-2)+in_buf[482]*(7)+in_buf[483]*(25)+in_buf[484]*(18)+in_buf[485]*(6)+in_buf[486]*(18)+in_buf[487]*(23)+in_buf[488]*(13)+in_buf[489]*(-13)+in_buf[490]*(-9)+in_buf[491]*(0)+in_buf[492]*(19)+in_buf[493]*(21)+in_buf[494]*(28)+in_buf[495]*(-3)+in_buf[496]*(4)+in_buf[497]*(2)+in_buf[498]*(-6)+in_buf[499]*(0)+in_buf[500]*(-25)+in_buf[501]*(16)+in_buf[502]*(-15)+in_buf[503]*(15)+in_buf[504]*(-3)+in_buf[505]*(-5)+in_buf[506]*(-18)+in_buf[507]*(1)+in_buf[508]*(3)+in_buf[509]*(-8)+in_buf[510]*(10)+in_buf[511]*(19)+in_buf[512]*(8)+in_buf[513]*(3)+in_buf[514]*(20)+in_buf[515]*(13)+in_buf[516]*(6)+in_buf[517]*(-5)+in_buf[518]*(-14)+in_buf[519]*(8)+in_buf[520]*(17)+in_buf[521]*(17)+in_buf[522]*(16)+in_buf[523]*(7)+in_buf[524]*(0)+in_buf[525]*(-2)+in_buf[526]*(-16)+in_buf[527]*(-9)+in_buf[528]*(-9)+in_buf[529]*(1)+in_buf[530]*(-28)+in_buf[531]*(-3)+in_buf[532]*(-5)+in_buf[533]*(-10)+in_buf[534]*(10)+in_buf[535]*(17)+in_buf[536]*(3)+in_buf[537]*(-1)+in_buf[538]*(0)+in_buf[539]*(7)+in_buf[540]*(9)+in_buf[541]*(-3)+in_buf[542]*(4)+in_buf[543]*(14)+in_buf[544]*(-4)+in_buf[545]*(-23)+in_buf[546]*(-2)+in_buf[547]*(13)+in_buf[548]*(16)+in_buf[549]*(0)+in_buf[550]*(16)+in_buf[551]*(6)+in_buf[552]*(-9)+in_buf[553]*(-7)+in_buf[554]*(-19)+in_buf[555]*(-8)+in_buf[556]*(12)+in_buf[557]*(4)+in_buf[558]*(14)+in_buf[559]*(7)+in_buf[560]*(-3)+in_buf[561]*(22)+in_buf[562]*(20)+in_buf[563]*(23)+in_buf[564]*(10)+in_buf[565]*(0)+in_buf[566]*(-9)+in_buf[567]*(-2)+in_buf[568]*(1)+in_buf[569]*(-15)+in_buf[570]*(3)+in_buf[571]*(-4)+in_buf[572]*(-15)+in_buf[573]*(-5)+in_buf[574]*(3)+in_buf[575]*(17)+in_buf[576]*(5)+in_buf[577]*(-4)+in_buf[578]*(5)+in_buf[579]*(-5)+in_buf[580]*(-15)+in_buf[581]*(-1)+in_buf[582]*(-12)+in_buf[583]*(-10)+in_buf[584]*(22)+in_buf[585]*(20)+in_buf[586]*(7)+in_buf[587]*(-2)+in_buf[588]*(-5)+in_buf[589]*(8)+in_buf[590]*(-13)+in_buf[591]*(11)+in_buf[592]*(23)+in_buf[593]*(16)+in_buf[594]*(1)+in_buf[595]*(4)+in_buf[596]*(2)+in_buf[597]*(1)+in_buf[598]*(-7)+in_buf[599]*(2)+in_buf[600]*(6)+in_buf[601]*(12)+in_buf[602]*(13)+in_buf[603]*(9)+in_buf[604]*(7)+in_buf[605]*(0)+in_buf[606]*(5)+in_buf[607]*(-2)+in_buf[608]*(-13)+in_buf[609]*(-9)+in_buf[610]*(-1)+in_buf[611]*(10)+in_buf[612]*(11)+in_buf[613]*(-9)+in_buf[614]*(15)+in_buf[615]*(0)+in_buf[616]*(0)+in_buf[617]*(1)+in_buf[618]*(-7)+in_buf[619]*(10)+in_buf[620]*(3)+in_buf[621]*(-21)+in_buf[622]*(-16)+in_buf[623]*(-4)+in_buf[624]*(-8)+in_buf[625]*(-12)+in_buf[626]*(-5)+in_buf[627]*(12)+in_buf[628]*(26)+in_buf[629]*(16)+in_buf[630]*(6)+in_buf[631]*(9)+in_buf[632]*(5)+in_buf[633]*(-12)+in_buf[634]*(-5)+in_buf[635]*(-5)+in_buf[636]*(-9)+in_buf[637]*(3)+in_buf[638]*(25)+in_buf[639]*(30)+in_buf[640]*(12)+in_buf[641]*(-13)+in_buf[642]*(3)+in_buf[643]*(1)+in_buf[644]*(0)+in_buf[645]*(1)+in_buf[646]*(-15)+in_buf[647]*(9)+in_buf[648]*(8)+in_buf[649]*(3)+in_buf[650]*(-7)+in_buf[651]*(-2)+in_buf[652]*(15)+in_buf[653]*(-6)+in_buf[654]*(-1)+in_buf[655]*(-2)+in_buf[656]*(-1)+in_buf[657]*(10)+in_buf[658]*(6)+in_buf[659]*(-6)+in_buf[660]*(-14)+in_buf[661]*(-17)+in_buf[662]*(-9)+in_buf[663]*(0)+in_buf[664]*(7)+in_buf[665]*(44)+in_buf[666]*(29)+in_buf[667]*(16)+in_buf[668]*(23)+in_buf[669]*(1)+in_buf[670]*(-5)+in_buf[671]*(-2)+in_buf[672]*(4)+in_buf[673]*(-3)+in_buf[674]*(-25)+in_buf[675]*(-20)+in_buf[676]*(-8)+in_buf[677]*(13)+in_buf[678]*(2)+in_buf[679]*(0)+in_buf[680]*(2)+in_buf[681]*(12)+in_buf[682]*(2)+in_buf[683]*(7)+in_buf[684]*(4)+in_buf[685]*(2)+in_buf[686]*(-4)+in_buf[687]*(0)+in_buf[688]*(-10)+in_buf[689]*(-13)+in_buf[690]*(-4)+in_buf[691]*(5)+in_buf[692]*(22)+in_buf[693]*(16)+in_buf[694]*(47)+in_buf[695]*(38)+in_buf[696]*(-11)+in_buf[697]*(14)+in_buf[698]*(-9)+in_buf[699]*(3)+in_buf[700]*(-1)+in_buf[701]*(-1)+in_buf[702]*(33)+in_buf[703]*(3)+in_buf[704]*(-9)+in_buf[705]*(6)+in_buf[706]*(6)+in_buf[707]*(-19)+in_buf[708]*(-13)+in_buf[709]*(-19)+in_buf[710]*(-13)+in_buf[711]*(-12)+in_buf[712]*(-28)+in_buf[713]*(-15)+in_buf[714]*(-5)+in_buf[715]*(-3)+in_buf[716]*(-23)+in_buf[717]*(-22)+in_buf[718]*(18)+in_buf[719]*(24)+in_buf[720]*(8)+in_buf[721]*(11)+in_buf[722]*(3)+in_buf[723]*(-13)+in_buf[724]*(-36)+in_buf[725]*(3)+in_buf[726]*(-9)+in_buf[727]*(-3)+in_buf[728]*(3)+in_buf[729]*(3)+in_buf[730]*(4)+in_buf[731]*(1)+in_buf[732]*(23)+in_buf[733]*(26)+in_buf[734]*(39)+in_buf[735]*(15)+in_buf[736]*(23)+in_buf[737]*(-3)+in_buf[738]*(3)+in_buf[739]*(-2)+in_buf[740]*(31)+in_buf[741]*(27)+in_buf[742]*(8)+in_buf[743]*(6)+in_buf[744]*(-7)+in_buf[745]*(-17)+in_buf[746]*(-6)+in_buf[747]*(-3)+in_buf[748]*(5)+in_buf[749]*(-3)+in_buf[750]*(6)+in_buf[751]*(30)+in_buf[752]*(20)+in_buf[753]*(0)+in_buf[754]*(3)+in_buf[755]*(-2)+in_buf[756]*(0)+in_buf[757]*(-1)+in_buf[758]*(-3)+in_buf[759]*(-2)+in_buf[760]*(-10)+in_buf[761]*(-12)+in_buf[762]*(-2)+in_buf[763]*(4)+in_buf[764]*(-1)+in_buf[765]*(-15)+in_buf[766]*(17)+in_buf[767]*(9)+in_buf[768]*(1)+in_buf[769]*(-33)+in_buf[770]*(-18)+in_buf[771]*(5)+in_buf[772]*(-19)+in_buf[773]*(-33)+in_buf[774]*(-17)+in_buf[775]*(26)+in_buf[776]*(26)+in_buf[777]*(0)+in_buf[778]*(-6)+in_buf[779]*(-26)+in_buf[780]*(3)+in_buf[781]*(0)+in_buf[782]*(1)+in_buf[783]*(4);
assign in_buf_weight025=in_buf[0]*(1)+in_buf[1]*(-3)+in_buf[2]*(0)+in_buf[3]*(2)+in_buf[4]*(2)+in_buf[5]*(1)+in_buf[6]*(4)+in_buf[7]*(1)+in_buf[8]*(-3)+in_buf[9]*(-1)+in_buf[10]*(0)+in_buf[11]*(-2)+in_buf[12]*(0)+in_buf[13]*(0)+in_buf[14]*(-2)+in_buf[15]*(0)+in_buf[16]*(3)+in_buf[17]*(1)+in_buf[18]*(0)+in_buf[19]*(-2)+in_buf[20]*(-3)+in_buf[21]*(-3)+in_buf[22]*(-1)+in_buf[23]*(0)+in_buf[24]*(-2)+in_buf[25]*(0)+in_buf[26]*(0)+in_buf[27]*(0)+in_buf[28]*(-2)+in_buf[29]*(0)+in_buf[30]*(4)+in_buf[31]*(1)+in_buf[32]*(1)+in_buf[33]*(-6)+in_buf[34]*(-12)+in_buf[35]*(-5)+in_buf[36]*(-11)+in_buf[37]*(-5)+in_buf[38]*(-8)+in_buf[39]*(-8)+in_buf[40]*(-16)+in_buf[41]*(-11)+in_buf[42]*(-6)+in_buf[43]*(-28)+in_buf[44]*(-27)+in_buf[45]*(-29)+in_buf[46]*(-10)+in_buf[47]*(-6)+in_buf[48]*(-8)+in_buf[49]*(-4)+in_buf[50]*(-3)+in_buf[51]*(-2)+in_buf[52]*(-3)+in_buf[53]*(1)+in_buf[54]*(0)+in_buf[55]*(-2)+in_buf[56]*(0)+in_buf[57]*(-1)+in_buf[58]*(-4)+in_buf[59]*(-1)+in_buf[60]*(-2)+in_buf[61]*(-2)+in_buf[62]*(-6)+in_buf[63]*(-11)+in_buf[64]*(-12)+in_buf[65]*(-21)+in_buf[66]*(-27)+in_buf[67]*(-13)+in_buf[68]*(-22)+in_buf[69]*(-35)+in_buf[70]*(-45)+in_buf[71]*(-19)+in_buf[72]*(-24)+in_buf[73]*(-4)+in_buf[74]*(-2)+in_buf[75]*(-8)+in_buf[76]*(-2)+in_buf[77]*(3)+in_buf[78]*(5)+in_buf[79]*(-22)+in_buf[80]*(-4)+in_buf[81]*(-1)+in_buf[82]*(5)+in_buf[83]*(4)+in_buf[84]*(-1)+in_buf[85]*(-1)+in_buf[86]*(2)+in_buf[87]*(-2)+in_buf[88]*(5)+in_buf[89]*(-21)+in_buf[90]*(-29)+in_buf[91]*(-36)+in_buf[92]*(-55)+in_buf[93]*(-44)+in_buf[94]*(-36)+in_buf[95]*(-33)+in_buf[96]*(-34)+in_buf[97]*(-50)+in_buf[98]*(-41)+in_buf[99]*(-1)+in_buf[100]*(23)+in_buf[101]*(6)+in_buf[102]*(16)+in_buf[103]*(39)+in_buf[104]*(24)+in_buf[105]*(2)+in_buf[106]*(-5)+in_buf[107]*(-9)+in_buf[108]*(-48)+in_buf[109]*(-28)+in_buf[110]*(-23)+in_buf[111]*(-4)+in_buf[112]*(3)+in_buf[113]*(4)+in_buf[114]*(0)+in_buf[115]*(31)+in_buf[116]*(27)+in_buf[117]*(28)+in_buf[118]*(-12)+in_buf[119]*(-7)+in_buf[120]*(-28)+in_buf[121]*(-33)+in_buf[122]*(4)+in_buf[123]*(15)+in_buf[124]*(25)+in_buf[125]*(4)+in_buf[126]*(-31)+in_buf[127]*(-23)+in_buf[128]*(1)+in_buf[129]*(-22)+in_buf[130]*(-13)+in_buf[131]*(22)+in_buf[132]*(2)+in_buf[133]*(6)+in_buf[134]*(6)+in_buf[135]*(-10)+in_buf[136]*(-3)+in_buf[137]*(-23)+in_buf[138]*(-3)+in_buf[139]*(-14)+in_buf[140]*(1)+in_buf[141]*(3)+in_buf[142]*(-15)+in_buf[143]*(4)+in_buf[144]*(-23)+in_buf[145]*(30)+in_buf[146]*(23)+in_buf[147]*(20)+in_buf[148]*(1)+in_buf[149]*(4)+in_buf[150]*(-21)+in_buf[151]*(0)+in_buf[152]*(10)+in_buf[153]*(-15)+in_buf[154]*(-12)+in_buf[155]*(-10)+in_buf[156]*(-14)+in_buf[157]*(-39)+in_buf[158]*(-19)+in_buf[159]*(0)+in_buf[160]*(5)+in_buf[161]*(7)+in_buf[162]*(7)+in_buf[163]*(-7)+in_buf[164]*(-6)+in_buf[165]*(2)+in_buf[166]*(-18)+in_buf[167]*(0)+in_buf[168]*(-2)+in_buf[169]*(-14)+in_buf[170]*(-10)+in_buf[171]*(-2)+in_buf[172]*(-3)+in_buf[173]*(20)+in_buf[174]*(26)+in_buf[175]*(11)+in_buf[176]*(8)+in_buf[177]*(0)+in_buf[178]*(-21)+in_buf[179]*(2)+in_buf[180]*(-7)+in_buf[181]*(-19)+in_buf[182]*(-20)+in_buf[183]*(-18)+in_buf[184]*(-15)+in_buf[185]*(-9)+in_buf[186]*(5)+in_buf[187]*(17)+in_buf[188]*(38)+in_buf[189]*(26)+in_buf[190]*(26)+in_buf[191]*(19)+in_buf[192]*(2)+in_buf[193]*(8)+in_buf[194]*(3)+in_buf[195]*(-21)+in_buf[196]*(2)+in_buf[197]*(-4)+in_buf[198]*(-4)+in_buf[199]*(23)+in_buf[200]*(2)+in_buf[201]*(-11)+in_buf[202]*(19)+in_buf[203]*(16)+in_buf[204]*(-2)+in_buf[205]*(0)+in_buf[206]*(5)+in_buf[207]*(-10)+in_buf[208]*(-11)+in_buf[209]*(-20)+in_buf[210]*(-33)+in_buf[211]*(-25)+in_buf[212]*(-7)+in_buf[213]*(14)+in_buf[214]*(18)+in_buf[215]*(22)+in_buf[216]*(38)+in_buf[217]*(21)+in_buf[218]*(17)+in_buf[219]*(22)+in_buf[220]*(7)+in_buf[221]*(-8)+in_buf[222]*(8)+in_buf[223]*(-20)+in_buf[224]*(-27)+in_buf[225]*(32)+in_buf[226]*(2)+in_buf[227]*(10)+in_buf[228]*(5)+in_buf[229]*(9)+in_buf[230]*(23)+in_buf[231]*(28)+in_buf[232]*(2)+in_buf[233]*(2)+in_buf[234]*(-3)+in_buf[235]*(-6)+in_buf[236]*(16)+in_buf[237]*(-3)+in_buf[238]*(-20)+in_buf[239]*(-12)+in_buf[240]*(-2)+in_buf[241]*(21)+in_buf[242]*(29)+in_buf[243]*(20)+in_buf[244]*(27)+in_buf[245]*(17)+in_buf[246]*(18)+in_buf[247]*(18)+in_buf[248]*(23)+in_buf[249]*(25)+in_buf[250]*(27)+in_buf[251]*(-3)+in_buf[252]*(16)+in_buf[253]*(26)+in_buf[254]*(0)+in_buf[255]*(5)+in_buf[256]*(23)+in_buf[257]*(13)+in_buf[258]*(21)+in_buf[259]*(17)+in_buf[260]*(12)+in_buf[261]*(2)+in_buf[262]*(-1)+in_buf[263]*(22)+in_buf[264]*(16)+in_buf[265]*(10)+in_buf[266]*(2)+in_buf[267]*(2)+in_buf[268]*(11)+in_buf[269]*(26)+in_buf[270]*(33)+in_buf[271]*(9)+in_buf[272]*(25)+in_buf[273]*(24)+in_buf[274]*(11)+in_buf[275]*(-9)+in_buf[276]*(2)+in_buf[277]*(14)+in_buf[278]*(13)+in_buf[279]*(-7)+in_buf[280]*(20)+in_buf[281]*(19)+in_buf[282]*(5)+in_buf[283]*(-18)+in_buf[284]*(30)+in_buf[285]*(2)+in_buf[286]*(0)+in_buf[287]*(10)+in_buf[288]*(6)+in_buf[289]*(17)+in_buf[290]*(20)+in_buf[291]*(30)+in_buf[292]*(24)+in_buf[293]*(-1)+in_buf[294]*(-14)+in_buf[295]*(0)+in_buf[296]*(3)+in_buf[297]*(18)+in_buf[298]*(11)+in_buf[299]*(2)+in_buf[300]*(-3)+in_buf[301]*(-9)+in_buf[302]*(-17)+in_buf[303]*(-43)+in_buf[304]*(-41)+in_buf[305]*(6)+in_buf[306]*(-31)+in_buf[307]*(7)+in_buf[308]*(20)+in_buf[309]*(-7)+in_buf[310]*(48)+in_buf[311]*(13)+in_buf[312]*(35)+in_buf[313]*(21)+in_buf[314]*(12)+in_buf[315]*(27)+in_buf[316]*(19)+in_buf[317]*(24)+in_buf[318]*(21)+in_buf[319]*(30)+in_buf[320]*(22)+in_buf[321]*(-13)+in_buf[322]*(-2)+in_buf[323]*(-7)+in_buf[324]*(1)+in_buf[325]*(1)+in_buf[326]*(2)+in_buf[327]*(-7)+in_buf[328]*(-6)+in_buf[329]*(-31)+in_buf[330]*(-31)+in_buf[331]*(-51)+in_buf[332]*(-58)+in_buf[333]*(-30)+in_buf[334]*(-41)+in_buf[335]*(25)+in_buf[336]*(21)+in_buf[337]*(21)+in_buf[338]*(22)+in_buf[339]*(35)+in_buf[340]*(35)+in_buf[341]*(25)+in_buf[342]*(9)+in_buf[343]*(30)+in_buf[344]*(24)+in_buf[345]*(4)+in_buf[346]*(10)+in_buf[347]*(18)+in_buf[348]*(3)+in_buf[349]*(2)+in_buf[350]*(5)+in_buf[351]*(14)+in_buf[352]*(13)+in_buf[353]*(7)+in_buf[354]*(5)+in_buf[355]*(-12)+in_buf[356]*(0)+in_buf[357]*(-16)+in_buf[358]*(-19)+in_buf[359]*(-34)+in_buf[360]*(-35)+in_buf[361]*(-22)+in_buf[362]*(-25)+in_buf[363]*(24)+in_buf[364]*(3)+in_buf[365]*(13)+in_buf[366]*(42)+in_buf[367]*(21)+in_buf[368]*(25)+in_buf[369]*(30)+in_buf[370]*(10)+in_buf[371]*(27)+in_buf[372]*(7)+in_buf[373]*(0)+in_buf[374]*(3)+in_buf[375]*(-1)+in_buf[376]*(-7)+in_buf[377]*(-3)+in_buf[378]*(14)+in_buf[379]*(30)+in_buf[380]*(20)+in_buf[381]*(9)+in_buf[382]*(2)+in_buf[383]*(-9)+in_buf[384]*(27)+in_buf[385]*(1)+in_buf[386]*(-15)+in_buf[387]*(-38)+in_buf[388]*(-26)+in_buf[389]*(-18)+in_buf[390]*(-38)+in_buf[391]*(-12)+in_buf[392]*(-3)+in_buf[393]*(15)+in_buf[394]*(39)+in_buf[395]*(13)+in_buf[396]*(19)+in_buf[397]*(24)+in_buf[398]*(-10)+in_buf[399]*(0)+in_buf[400]*(-11)+in_buf[401]*(-4)+in_buf[402]*(5)+in_buf[403]*(-7)+in_buf[404]*(-8)+in_buf[405]*(-5)+in_buf[406]*(15)+in_buf[407]*(7)+in_buf[408]*(17)+in_buf[409]*(6)+in_buf[410]*(-3)+in_buf[411]*(20)+in_buf[412]*(5)+in_buf[413]*(-10)+in_buf[414]*(1)+in_buf[415]*(14)+in_buf[416]*(-19)+in_buf[417]*(-46)+in_buf[418]*(-52)+in_buf[419]*(-17)+in_buf[420]*(5)+in_buf[421]*(7)+in_buf[422]*(29)+in_buf[423]*(34)+in_buf[424]*(0)+in_buf[425]*(-13)+in_buf[426]*(-6)+in_buf[427]*(4)+in_buf[428]*(-4)+in_buf[429]*(10)+in_buf[430]*(15)+in_buf[431]*(0)+in_buf[432]*(-24)+in_buf[433]*(-7)+in_buf[434]*(17)+in_buf[435]*(15)+in_buf[436]*(9)+in_buf[437]*(12)+in_buf[438]*(9)+in_buf[439]*(15)+in_buf[440]*(11)+in_buf[441]*(-2)+in_buf[442]*(37)+in_buf[443]*(28)+in_buf[444]*(-28)+in_buf[445]*(-38)+in_buf[446]*(-10)+in_buf[447]*(-2)+in_buf[448]*(10)+in_buf[449]*(0)+in_buf[450]*(20)+in_buf[451]*(6)+in_buf[452]*(-20)+in_buf[453]*(-24)+in_buf[454]*(13)+in_buf[455]*(13)+in_buf[456]*(-3)+in_buf[457]*(19)+in_buf[458]*(6)+in_buf[459]*(-19)+in_buf[460]*(0)+in_buf[461]*(5)+in_buf[462]*(22)+in_buf[463]*(12)+in_buf[464]*(15)+in_buf[465]*(23)+in_buf[466]*(12)+in_buf[467]*(5)+in_buf[468]*(14)+in_buf[469]*(18)+in_buf[470]*(8)+in_buf[471]*(-2)+in_buf[472]*(-18)+in_buf[473]*(-36)+in_buf[474]*(-49)+in_buf[475]*(-23)+in_buf[476]*(2)+in_buf[477]*(10)+in_buf[478]*(14)+in_buf[479]*(-21)+in_buf[480]*(-12)+in_buf[481]*(-21)+in_buf[482]*(0)+in_buf[483]*(-2)+in_buf[484]*(-2)+in_buf[485]*(-2)+in_buf[486]*(-9)+in_buf[487]*(-14)+in_buf[488]*(-11)+in_buf[489]*(-8)+in_buf[490]*(15)+in_buf[491]*(16)+in_buf[492]*(11)+in_buf[493]*(17)+in_buf[494]*(0)+in_buf[495]*(-18)+in_buf[496]*(3)+in_buf[497]*(15)+in_buf[498]*(3)+in_buf[499]*(-6)+in_buf[500]*(3)+in_buf[501]*(-17)+in_buf[502]*(-48)+in_buf[503]*(-19)+in_buf[504]*(32)+in_buf[505]*(3)+in_buf[506]*(31)+in_buf[507]*(-14)+in_buf[508]*(-7)+in_buf[509]*(-19)+in_buf[510]*(-17)+in_buf[511]*(-10)+in_buf[512]*(-11)+in_buf[513]*(-17)+in_buf[514]*(-36)+in_buf[515]*(-28)+in_buf[516]*(-19)+in_buf[517]*(-2)+in_buf[518]*(4)+in_buf[519]*(9)+in_buf[520]*(5)+in_buf[521]*(-2)+in_buf[522]*(-20)+in_buf[523]*(-9)+in_buf[524]*(4)+in_buf[525]*(5)+in_buf[526]*(-6)+in_buf[527]*(-17)+in_buf[528]*(-20)+in_buf[529]*(-14)+in_buf[530]*(5)+in_buf[531]*(8)+in_buf[532]*(9)+in_buf[533]*(32)+in_buf[534]*(24)+in_buf[535]*(-18)+in_buf[536]*(-7)+in_buf[537]*(-31)+in_buf[538]*(-29)+in_buf[539]*(-19)+in_buf[540]*(-2)+in_buf[541]*(-19)+in_buf[542]*(-49)+in_buf[543]*(-47)+in_buf[544]*(-37)+in_buf[545]*(-14)+in_buf[546]*(4)+in_buf[547]*(5)+in_buf[548]*(3)+in_buf[549]*(0)+in_buf[550]*(-18)+in_buf[551]*(8)+in_buf[552]*(-8)+in_buf[553]*(-9)+in_buf[554]*(-15)+in_buf[555]*(-23)+in_buf[556]*(-36)+in_buf[557]*(-31)+in_buf[558]*(-7)+in_buf[559]*(16)+in_buf[560]*(0)+in_buf[561]*(0)+in_buf[562]*(1)+in_buf[563]*(-41)+in_buf[564]*(-47)+in_buf[565]*(-42)+in_buf[566]*(-21)+in_buf[567]*(-17)+in_buf[568]*(-3)+in_buf[569]*(-25)+in_buf[570]*(-26)+in_buf[571]*(-42)+in_buf[572]*(-36)+in_buf[573]*(-20)+in_buf[574]*(1)+in_buf[575]*(13)+in_buf[576]*(8)+in_buf[577]*(10)+in_buf[578]*(0)+in_buf[579]*(-3)+in_buf[580]*(-11)+in_buf[581]*(-12)+in_buf[582]*(-4)+in_buf[583]*(-16)+in_buf[584]*(-26)+in_buf[585]*(-38)+in_buf[586]*(-11)+in_buf[587]*(8)+in_buf[588]*(7)+in_buf[589]*(3)+in_buf[590]*(1)+in_buf[591]*(-34)+in_buf[592]*(-20)+in_buf[593]*(-1)+in_buf[594]*(2)+in_buf[595]*(3)+in_buf[596]*(1)+in_buf[597]*(-3)+in_buf[598]*(-10)+in_buf[599]*(-12)+in_buf[600]*(-9)+in_buf[601]*(-4)+in_buf[602]*(2)+in_buf[603]*(18)+in_buf[604]*(0)+in_buf[605]*(11)+in_buf[606]*(0)+in_buf[607]*(-4)+in_buf[608]*(9)+in_buf[609]*(12)+in_buf[610]*(-1)+in_buf[611]*(-11)+in_buf[612]*(-13)+in_buf[613]*(12)+in_buf[614]*(-25)+in_buf[615]*(2)+in_buf[616]*(2)+in_buf[617]*(7)+in_buf[618]*(-14)+in_buf[619]*(-45)+in_buf[620]*(3)+in_buf[621]*(26)+in_buf[622]*(6)+in_buf[623]*(3)+in_buf[624]*(0)+in_buf[625]*(1)+in_buf[626]*(0)+in_buf[627]*(2)+in_buf[628]*(0)+in_buf[629]*(4)+in_buf[630]*(15)+in_buf[631]*(18)+in_buf[632]*(12)+in_buf[633]*(10)+in_buf[634]*(9)+in_buf[635]*(31)+in_buf[636]*(21)+in_buf[637]*(7)+in_buf[638]*(-11)+in_buf[639]*(-17)+in_buf[640]*(-15)+in_buf[641]*(8)+in_buf[642]*(4)+in_buf[643]*(-5)+in_buf[644]*(0)+in_buf[645]*(0)+in_buf[646]*(-18)+in_buf[647]*(-48)+in_buf[648]*(8)+in_buf[649]*(9)+in_buf[650]*(8)+in_buf[651]*(11)+in_buf[652]*(-11)+in_buf[653]*(2)+in_buf[654]*(7)+in_buf[655]*(-3)+in_buf[656]*(-2)+in_buf[657]*(0)+in_buf[658]*(6)+in_buf[659]*(17)+in_buf[660]*(16)+in_buf[661]*(5)+in_buf[662]*(11)+in_buf[663]*(23)+in_buf[664]*(-9)+in_buf[665]*(-19)+in_buf[666]*(-22)+in_buf[667]*(-21)+in_buf[668]*(-37)+in_buf[669]*(-30)+in_buf[670]*(27)+in_buf[671]*(0)+in_buf[672]*(-3)+in_buf[673]*(-2)+in_buf[674]*(5)+in_buf[675]*(-16)+in_buf[676]*(9)+in_buf[677]*(16)+in_buf[678]*(6)+in_buf[679]*(2)+in_buf[680]*(-4)+in_buf[681]*(-5)+in_buf[682]*(11)+in_buf[683]*(17)+in_buf[684]*(1)+in_buf[685]*(10)+in_buf[686]*(9)+in_buf[687]*(13)+in_buf[688]*(2)+in_buf[689]*(-17)+in_buf[690]*(-12)+in_buf[691]*(0)+in_buf[692]*(-7)+in_buf[693]*(-21)+in_buf[694]*(-20)+in_buf[695]*(-19)+in_buf[696]*(-26)+in_buf[697]*(-24)+in_buf[698]*(-7)+in_buf[699]*(-1)+in_buf[700]*(0)+in_buf[701]*(-2)+in_buf[702]*(-24)+in_buf[703]*(11)+in_buf[704]*(28)+in_buf[705]*(0)+in_buf[706]*(-1)+in_buf[707]*(1)+in_buf[708]*(28)+in_buf[709]*(22)+in_buf[710]*(-4)+in_buf[711]*(0)+in_buf[712]*(20)+in_buf[713]*(10)+in_buf[714]*(19)+in_buf[715]*(9)+in_buf[716]*(-5)+in_buf[717]*(-9)+in_buf[718]*(-5)+in_buf[719]*(-19)+in_buf[720]*(-9)+in_buf[721]*(2)+in_buf[722]*(1)+in_buf[723]*(-8)+in_buf[724]*(-28)+in_buf[725]*(-11)+in_buf[726]*(-4)+in_buf[727]*(-3)+in_buf[728]*(0)+in_buf[729]*(-2)+in_buf[730]*(1)+in_buf[731]*(-14)+in_buf[732]*(-37)+in_buf[733]*(-36)+in_buf[734]*(2)+in_buf[735]*(20)+in_buf[736]*(16)+in_buf[737]*(34)+in_buf[738]*(15)+in_buf[739]*(0)+in_buf[740]*(-8)+in_buf[741]*(0)+in_buf[742]*(18)+in_buf[743]*(23)+in_buf[744]*(-3)+in_buf[745]*(0)+in_buf[746]*(2)+in_buf[747]*(9)+in_buf[748]*(7)+in_buf[749]*(3)+in_buf[750]*(-11)+in_buf[751]*(3)+in_buf[752]*(0)+in_buf[753]*(11)+in_buf[754]*(0)+in_buf[755]*(2)+in_buf[756]*(2)+in_buf[757]*(-1)+in_buf[758]*(2)+in_buf[759]*(2)+in_buf[760]*(29)+in_buf[761]*(22)+in_buf[762]*(6)+in_buf[763]*(-4)+in_buf[764]*(-1)+in_buf[765]*(28)+in_buf[766]*(23)+in_buf[767]*(21)+in_buf[768]*(11)+in_buf[769]*(50)+in_buf[770]*(22)+in_buf[771]*(13)+in_buf[772]*(26)+in_buf[773]*(50)+in_buf[774]*(19)+in_buf[775]*(3)+in_buf[776]*(-2)+in_buf[777]*(22)+in_buf[778]*(7)+in_buf[779]*(32)+in_buf[780]*(2)+in_buf[781]*(2)+in_buf[782]*(4)+in_buf[783]*(0);
assign in_buf_weight026=in_buf[0]*(-1)+in_buf[1]*(-1)+in_buf[2]*(-3)+in_buf[3]*(-3)+in_buf[4]*(-1)+in_buf[5]*(-3)+in_buf[6]*(0)+in_buf[7]*(2)+in_buf[8]*(2)+in_buf[9]*(-3)+in_buf[10]*(4)+in_buf[11]*(-3)+in_buf[12]*(-3)+in_buf[13]*(9)+in_buf[14]*(19)+in_buf[15]*(16)+in_buf[16]*(2)+in_buf[17]*(0)+in_buf[18]*(-2)+in_buf[19]*(4)+in_buf[20]*(-1)+in_buf[21]*(4)+in_buf[22]*(2)+in_buf[23]*(-3)+in_buf[24]*(3)+in_buf[25]*(-3)+in_buf[26]*(-2)+in_buf[27]*(-3)+in_buf[28]*(0)+in_buf[29]*(0)+in_buf[30]*(-3)+in_buf[31]*(-1)+in_buf[32]*(1)+in_buf[33]*(3)+in_buf[34]*(13)+in_buf[35]*(6)+in_buf[36]*(5)+in_buf[37]*(4)+in_buf[38]*(4)+in_buf[39]*(9)+in_buf[40]*(12)+in_buf[41]*(-10)+in_buf[42]*(-11)+in_buf[43]*(23)+in_buf[44]*(8)+in_buf[45]*(19)+in_buf[46]*(-3)+in_buf[47]*(2)+in_buf[48]*(11)+in_buf[49]*(1)+in_buf[50]*(3)+in_buf[51]*(6)+in_buf[52]*(-1)+in_buf[53]*(3)+in_buf[54]*(-2)+in_buf[55]*(1)+in_buf[56]*(-2)+in_buf[57]*(2)+in_buf[58]*(16)+in_buf[59]*(0)+in_buf[60]*(12)+in_buf[61]*(7)+in_buf[62]*(4)+in_buf[63]*(5)+in_buf[64]*(7)+in_buf[65]*(32)+in_buf[66]*(45)+in_buf[67]*(24)+in_buf[68]*(13)+in_buf[69]*(-1)+in_buf[70]*(-9)+in_buf[71]*(17)+in_buf[72]*(45)+in_buf[73]*(36)+in_buf[74]*(2)+in_buf[75]*(26)+in_buf[76]*(24)+in_buf[77]*(13)+in_buf[78]*(-4)+in_buf[79]*(33)+in_buf[80]*(10)+in_buf[81]*(12)+in_buf[82]*(0)+in_buf[83]*(3)+in_buf[84]*(-2)+in_buf[85]*(2)+in_buf[86]*(29)+in_buf[87]*(16)+in_buf[88]*(27)+in_buf[89]*(2)+in_buf[90]*(0)+in_buf[91]*(1)+in_buf[92]*(38)+in_buf[93]*(33)+in_buf[94]*(9)+in_buf[95]*(12)+in_buf[96]*(18)+in_buf[97]*(0)+in_buf[98]*(-39)+in_buf[99]*(-33)+in_buf[100]*(-10)+in_buf[101]*(-6)+in_buf[102]*(12)+in_buf[103]*(22)+in_buf[104]*(5)+in_buf[105]*(-2)+in_buf[106]*(1)+in_buf[107]*(-22)+in_buf[108]*(10)+in_buf[109]*(22)+in_buf[110]*(9)+in_buf[111]*(0)+in_buf[112]*(4)+in_buf[113]*(7)+in_buf[114]*(28)+in_buf[115]*(32)+in_buf[116]*(-2)+in_buf[117]*(16)+in_buf[118]*(5)+in_buf[119]*(-11)+in_buf[120]*(17)+in_buf[121]*(-14)+in_buf[122]*(-5)+in_buf[123]*(10)+in_buf[124]*(4)+in_buf[125]*(3)+in_buf[126]*(12)+in_buf[127]*(5)+in_buf[128]*(1)+in_buf[129]*(-10)+in_buf[130]*(1)+in_buf[131]*(23)+in_buf[132]*(0)+in_buf[133]*(-13)+in_buf[134]*(-1)+in_buf[135]*(0)+in_buf[136]*(-7)+in_buf[137]*(27)+in_buf[138]*(4)+in_buf[139]*(-13)+in_buf[140]*(0)+in_buf[141]*(0)+in_buf[142]*(18)+in_buf[143]*(3)+in_buf[144]*(4)+in_buf[145]*(17)+in_buf[146]*(8)+in_buf[147]*(-4)+in_buf[148]*(-2)+in_buf[149]*(-7)+in_buf[150]*(-16)+in_buf[151]*(-13)+in_buf[152]*(-16)+in_buf[153]*(-15)+in_buf[154]*(-7)+in_buf[155]*(0)+in_buf[156]*(2)+in_buf[157]*(-15)+in_buf[158]*(-14)+in_buf[159]*(5)+in_buf[160]*(18)+in_buf[161]*(10)+in_buf[162]*(20)+in_buf[163]*(29)+in_buf[164]*(7)+in_buf[165]*(2)+in_buf[166]*(17)+in_buf[167]*(-9)+in_buf[168]*(0)+in_buf[169]*(25)+in_buf[170]*(-7)+in_buf[171]*(-9)+in_buf[172]*(9)+in_buf[173]*(18)+in_buf[174]*(25)+in_buf[175]*(28)+in_buf[176]*(22)+in_buf[177]*(17)+in_buf[178]*(12)+in_buf[179]*(9)+in_buf[180]*(-1)+in_buf[181]*(-10)+in_buf[182]*(-15)+in_buf[183]*(-6)+in_buf[184]*(-11)+in_buf[185]*(-21)+in_buf[186]*(-11)+in_buf[187]*(-1)+in_buf[188]*(-1)+in_buf[189]*(-4)+in_buf[190]*(12)+in_buf[191]*(20)+in_buf[192]*(31)+in_buf[193]*(23)+in_buf[194]*(41)+in_buf[195]*(36)+in_buf[196]*(0)+in_buf[197]*(47)+in_buf[198]*(-4)+in_buf[199]*(3)+in_buf[200]*(28)+in_buf[201]*(23)+in_buf[202]*(20)+in_buf[203]*(29)+in_buf[204]*(23)+in_buf[205]*(19)+in_buf[206]*(22)+in_buf[207]*(9)+in_buf[208]*(15)+in_buf[209]*(12)+in_buf[210]*(-2)+in_buf[211]*(-20)+in_buf[212]*(-8)+in_buf[213]*(-1)+in_buf[214]*(8)+in_buf[215]*(13)+in_buf[216]*(16)+in_buf[217]*(8)+in_buf[218]*(9)+in_buf[219]*(6)+in_buf[220]*(2)+in_buf[221]*(24)+in_buf[222]*(60)+in_buf[223]*(33)+in_buf[224]*(-1)+in_buf[225]*(28)+in_buf[226]*(-9)+in_buf[227]*(12)+in_buf[228]*(17)+in_buf[229]*(8)+in_buf[230]*(-11)+in_buf[231]*(21)+in_buf[232]*(5)+in_buf[233]*(19)+in_buf[234]*(21)+in_buf[235]*(28)+in_buf[236]*(25)+in_buf[237]*(11)+in_buf[238]*(-4)+in_buf[239]*(-12)+in_buf[240]*(-9)+in_buf[241]*(17)+in_buf[242]*(4)+in_buf[243]*(23)+in_buf[244]*(29)+in_buf[245]*(1)+in_buf[246]*(25)+in_buf[247]*(28)+in_buf[248]*(0)+in_buf[249]*(11)+in_buf[250]*(49)+in_buf[251]*(10)+in_buf[252]*(-2)+in_buf[253]*(21)+in_buf[254]*(3)+in_buf[255]*(18)+in_buf[256]*(11)+in_buf[257]*(0)+in_buf[258]*(-11)+in_buf[259]*(19)+in_buf[260]*(17)+in_buf[261]*(2)+in_buf[262]*(1)+in_buf[263]*(16)+in_buf[264]*(13)+in_buf[265]*(-18)+in_buf[266]*(-21)+in_buf[267]*(-11)+in_buf[268]*(8)+in_buf[269]*(14)+in_buf[270]*(15)+in_buf[271]*(12)+in_buf[272]*(3)+in_buf[273]*(8)+in_buf[274]*(43)+in_buf[275]*(20)+in_buf[276]*(0)+in_buf[277]*(3)+in_buf[278]*(47)+in_buf[279]*(32)+in_buf[280]*(-1)+in_buf[281]*(24)+in_buf[282]*(2)+in_buf[283]*(-4)+in_buf[284]*(-2)+in_buf[285]*(-25)+in_buf[286]*(-6)+in_buf[287]*(7)+in_buf[288]*(12)+in_buf[289]*(-7)+in_buf[290]*(-4)+in_buf[291]*(-12)+in_buf[292]*(-30)+in_buf[293]*(-44)+in_buf[294]*(-32)+in_buf[295]*(-19)+in_buf[296]*(6)+in_buf[297]*(8)+in_buf[298]*(7)+in_buf[299]*(-5)+in_buf[300]*(-7)+in_buf[301]*(8)+in_buf[302]*(16)+in_buf[303]*(-6)+in_buf[304]*(6)+in_buf[305]*(18)+in_buf[306]*(28)+in_buf[307]*(28)+in_buf[308]*(-1)+in_buf[309]*(21)+in_buf[310]*(-22)+in_buf[311]*(-21)+in_buf[312]*(-20)+in_buf[313]*(-25)+in_buf[314]*(-40)+in_buf[315]*(-16)+in_buf[316]*(-31)+in_buf[317]*(-44)+in_buf[318]*(-53)+in_buf[319]*(-32)+in_buf[320]*(-63)+in_buf[321]*(-39)+in_buf[322]*(1)+in_buf[323]*(-2)+in_buf[324]*(-7)+in_buf[325]*(-6)+in_buf[326]*(-12)+in_buf[327]*(-23)+in_buf[328]*(-27)+in_buf[329]*(-10)+in_buf[330]*(-6)+in_buf[331]*(-12)+in_buf[332]*(8)+in_buf[333]*(24)+in_buf[334]*(-1)+in_buf[335]*(37)+in_buf[336]*(-1)+in_buf[337]*(-11)+in_buf[338]*(-32)+in_buf[339]*(-30)+in_buf[340]*(-47)+in_buf[341]*(-63)+in_buf[342]*(-78)+in_buf[343]*(-63)+in_buf[344]*(-68)+in_buf[345]*(-81)+in_buf[346]*(-59)+in_buf[347]*(-49)+in_buf[348]*(-34)+in_buf[349]*(-7)+in_buf[350]*(21)+in_buf[351]*(4)+in_buf[352]*(-1)+in_buf[353]*(-17)+in_buf[354]*(-15)+in_buf[355]*(-20)+in_buf[356]*(-15)+in_buf[357]*(-8)+in_buf[358]*(-20)+in_buf[359]*(-23)+in_buf[360]*(-1)+in_buf[361]*(18)+in_buf[362]*(8)+in_buf[363]*(34)+in_buf[364]*(5)+in_buf[365]*(-17)+in_buf[366]*(-18)+in_buf[367]*(-33)+in_buf[368]*(-72)+in_buf[369]*(-68)+in_buf[370]*(-69)+in_buf[371]*(-76)+in_buf[372]*(-57)+in_buf[373]*(-46)+in_buf[374]*(-38)+in_buf[375]*(-24)+in_buf[376]*(12)+in_buf[377]*(29)+in_buf[378]*(26)+in_buf[379]*(8)+in_buf[380]*(7)+in_buf[381]*(-3)+in_buf[382]*(-20)+in_buf[383]*(-10)+in_buf[384]*(0)+in_buf[385]*(2)+in_buf[386]*(-6)+in_buf[387]*(-15)+in_buf[388]*(-1)+in_buf[389]*(2)+in_buf[390]*(15)+in_buf[391]*(14)+in_buf[392]*(4)+in_buf[393]*(-17)+in_buf[394]*(-8)+in_buf[395]*(-27)+in_buf[396]*(-45)+in_buf[397]*(-32)+in_buf[398]*(-14)+in_buf[399]*(-22)+in_buf[400]*(-11)+in_buf[401]*(-7)+in_buf[402]*(7)+in_buf[403]*(18)+in_buf[404]*(36)+in_buf[405]*(41)+in_buf[406]*(29)+in_buf[407]*(2)+in_buf[408]*(6)+in_buf[409]*(3)+in_buf[410]*(2)+in_buf[411]*(13)+in_buf[412]*(-4)+in_buf[413]*(-3)+in_buf[414]*(5)+in_buf[415]*(-9)+in_buf[416]*(7)+in_buf[417]*(-12)+in_buf[418]*(34)+in_buf[419]*(12)+in_buf[420]*(4)+in_buf[421]*(4)+in_buf[422]*(19)+in_buf[423]*(-9)+in_buf[424]*(3)+in_buf[425]*(22)+in_buf[426]*(23)+in_buf[427]*(12)+in_buf[428]*(9)+in_buf[429]*(13)+in_buf[430]*(18)+in_buf[431]*(29)+in_buf[432]*(30)+in_buf[433]*(41)+in_buf[434]*(22)+in_buf[435]*(1)+in_buf[436]*(-6)+in_buf[437]*(5)+in_buf[438]*(18)+in_buf[439]*(7)+in_buf[440]*(-9)+in_buf[441]*(-2)+in_buf[442]*(-4)+in_buf[443]*(9)+in_buf[444]*(31)+in_buf[445]*(-7)+in_buf[446]*(-11)+in_buf[447]*(12)+in_buf[448]*(3)+in_buf[449]*(17)+in_buf[450]*(38)+in_buf[451]*(21)+in_buf[452]*(27)+in_buf[453]*(35)+in_buf[454]*(35)+in_buf[455]*(18)+in_buf[456]*(14)+in_buf[457]*(30)+in_buf[458]*(23)+in_buf[459]*(24)+in_buf[460]*(27)+in_buf[461]*(28)+in_buf[462]*(19)+in_buf[463]*(-4)+in_buf[464]*(-2)+in_buf[465]*(-3)+in_buf[466]*(8)+in_buf[467]*(18)+in_buf[468]*(-10)+in_buf[469]*(8)+in_buf[470]*(14)+in_buf[471]*(15)+in_buf[472]*(37)+in_buf[473]*(0)+in_buf[474]*(10)+in_buf[475]*(19)+in_buf[476]*(0)+in_buf[477]*(5)+in_buf[478]*(29)+in_buf[479]*(33)+in_buf[480]*(11)+in_buf[481]*(13)+in_buf[482]*(33)+in_buf[483]*(17)+in_buf[484]*(20)+in_buf[485]*(17)+in_buf[486]*(26)+in_buf[487]*(21)+in_buf[488]*(14)+in_buf[489]*(10)+in_buf[490]*(9)+in_buf[491]*(-10)+in_buf[492]*(-2)+in_buf[493]*(-9)+in_buf[494]*(5)+in_buf[495]*(11)+in_buf[496]*(-8)+in_buf[497]*(10)+in_buf[498]*(18)+in_buf[499]*(3)+in_buf[500]*(9)+in_buf[501]*(4)+in_buf[502]*(11)+in_buf[503]*(8)+in_buf[504]*(1)+in_buf[505]*(12)+in_buf[506]*(4)+in_buf[507]*(46)+in_buf[508]*(3)+in_buf[509]*(10)+in_buf[510]*(19)+in_buf[511]*(29)+in_buf[512]*(26)+in_buf[513]*(23)+in_buf[514]*(17)+in_buf[515]*(3)+in_buf[516]*(6)+in_buf[517]*(5)+in_buf[518]*(1)+in_buf[519]*(-5)+in_buf[520]*(1)+in_buf[521]*(5)+in_buf[522]*(5)+in_buf[523]*(0)+in_buf[524]*(-2)+in_buf[525]*(-4)+in_buf[526]*(3)+in_buf[527]*(-4)+in_buf[528]*(34)+in_buf[529]*(55)+in_buf[530]*(46)+in_buf[531]*(23)+in_buf[532]*(18)+in_buf[533]*(-27)+in_buf[534]*(-21)+in_buf[535]*(7)+in_buf[536]*(-4)+in_buf[537]*(-5)+in_buf[538]*(11)+in_buf[539]*(19)+in_buf[540]*(13)+in_buf[541]*(15)+in_buf[542]*(11)+in_buf[543]*(8)+in_buf[544]*(-3)+in_buf[545]*(7)+in_buf[546]*(6)+in_buf[547]*(-6)+in_buf[548]*(-5)+in_buf[549]*(11)+in_buf[550]*(4)+in_buf[551]*(9)+in_buf[552]*(-2)+in_buf[553]*(-7)+in_buf[554]*(-3)+in_buf[555]*(8)+in_buf[556]*(14)+in_buf[557]*(56)+in_buf[558]*(-5)+in_buf[559]*(16)+in_buf[560]*(-2)+in_buf[561]*(-30)+in_buf[562]*(-3)+in_buf[563]*(12)+in_buf[564]*(-9)+in_buf[565]*(-8)+in_buf[566]*(20)+in_buf[567]*(26)+in_buf[568]*(15)+in_buf[569]*(5)+in_buf[570]*(7)+in_buf[571]*(-2)+in_buf[572]*(3)+in_buf[573]*(9)+in_buf[574]*(9)+in_buf[575]*(-3)+in_buf[576]*(9)+in_buf[577]*(11)+in_buf[578]*(16)+in_buf[579]*(0)+in_buf[580]*(1)+in_buf[581]*(-7)+in_buf[582]*(-16)+in_buf[583]*(-1)+in_buf[584]*(-1)+in_buf[585]*(24)+in_buf[586]*(-4)+in_buf[587]*(2)+in_buf[588]*(24)+in_buf[589]*(17)+in_buf[590]*(35)+in_buf[591]*(33)+in_buf[592]*(-11)+in_buf[593]*(-2)+in_buf[594]*(0)+in_buf[595]*(14)+in_buf[596]*(3)+in_buf[597]*(-1)+in_buf[598]*(5)+in_buf[599]*(0)+in_buf[600]*(7)+in_buf[601]*(4)+in_buf[602]*(6)+in_buf[603]*(7)+in_buf[604]*(9)+in_buf[605]*(10)+in_buf[606]*(7)+in_buf[607]*(5)+in_buf[608]*(3)+in_buf[609]*(-6)+in_buf[610]*(-21)+in_buf[611]*(-7)+in_buf[612]*(4)+in_buf[613]*(27)+in_buf[614]*(27)+in_buf[615]*(0)+in_buf[616]*(21)+in_buf[617]*(19)+in_buf[618]*(49)+in_buf[619]*(26)+in_buf[620]*(12)+in_buf[621]*(17)+in_buf[622]*(-6)+in_buf[623]*(-1)+in_buf[624]*(-6)+in_buf[625]*(0)+in_buf[626]*(-2)+in_buf[627]*(-4)+in_buf[628]*(3)+in_buf[629]*(10)+in_buf[630]*(2)+in_buf[631]*(-1)+in_buf[632]*(5)+in_buf[633]*(10)+in_buf[634]*(1)+in_buf[635]*(18)+in_buf[636]*(17)+in_buf[637]*(-7)+in_buf[638]*(-20)+in_buf[639]*(-10)+in_buf[640]*(2)+in_buf[641]*(11)+in_buf[642]*(15)+in_buf[643]*(-5)+in_buf[644]*(2)+in_buf[645]*(-4)+in_buf[646]*(43)+in_buf[647]*(5)+in_buf[648]*(19)+in_buf[649]*(11)+in_buf[650]*(5)+in_buf[651]*(0)+in_buf[652]*(-10)+in_buf[653]*(0)+in_buf[654]*(-8)+in_buf[655]*(7)+in_buf[656]*(20)+in_buf[657]*(24)+in_buf[658]*(9)+in_buf[659]*(0)+in_buf[660]*(5)+in_buf[661]*(-4)+in_buf[662]*(-15)+in_buf[663]*(-14)+in_buf[664]*(-8)+in_buf[665]*(-3)+in_buf[666]*(9)+in_buf[667]*(13)+in_buf[668]*(12)+in_buf[669]*(18)+in_buf[670]*(30)+in_buf[671]*(-1)+in_buf[672]*(4)+in_buf[673]*(-1)+in_buf[674]*(26)+in_buf[675]*(5)+in_buf[676]*(17)+in_buf[677]*(-12)+in_buf[678]*(-12)+in_buf[679]*(-4)+in_buf[680]*(-3)+in_buf[681]*(5)+in_buf[682]*(-11)+in_buf[683]*(10)+in_buf[684]*(20)+in_buf[685]*(9)+in_buf[686]*(9)+in_buf[687]*(-20)+in_buf[688]*(0)+in_buf[689]*(-8)+in_buf[690]*(-22)+in_buf[691]*(-26)+in_buf[692]*(-2)+in_buf[693]*(-21)+in_buf[694]*(-23)+in_buf[695]*(-22)+in_buf[696]*(18)+in_buf[697]*(0)+in_buf[698]*(11)+in_buf[699]*(0)+in_buf[700]*(4)+in_buf[701]*(4)+in_buf[702]*(-21)+in_buf[703]*(16)+in_buf[704]*(6)+in_buf[705]*(-15)+in_buf[706]*(-6)+in_buf[707]*(2)+in_buf[708]*(9)+in_buf[709]*(17)+in_buf[710]*(14)+in_buf[711]*(5)+in_buf[712]*(26)+in_buf[713]*(5)+in_buf[714]*(0)+in_buf[715]*(2)+in_buf[716]*(5)+in_buf[717]*(3)+in_buf[718]*(-30)+in_buf[719]*(-32)+in_buf[720]*(-19)+in_buf[721]*(-54)+in_buf[722]*(-50)+in_buf[723]*(-11)+in_buf[724]*(3)+in_buf[725]*(-2)+in_buf[726]*(6)+in_buf[727]*(-3)+in_buf[728]*(3)+in_buf[729]*(-1)+in_buf[730]*(2)+in_buf[731]*(-1)+in_buf[732]*(-8)+in_buf[733]*(-26)+in_buf[734]*(-37)+in_buf[735]*(-5)+in_buf[736]*(-35)+in_buf[737]*(5)+in_buf[738]*(0)+in_buf[739]*(-4)+in_buf[740]*(-22)+in_buf[741]*(-12)+in_buf[742]*(-30)+in_buf[743]*(-27)+in_buf[744]*(-35)+in_buf[745]*(-14)+in_buf[746]*(-26)+in_buf[747]*(-8)+in_buf[748]*(-13)+in_buf[749]*(-25)+in_buf[750]*(-23)+in_buf[751]*(0)+in_buf[752]*(-1)+in_buf[753]*(3)+in_buf[754]*(4)+in_buf[755]*(3)+in_buf[756]*(4)+in_buf[757]*(0)+in_buf[758]*(2)+in_buf[759]*(-1)+in_buf[760]*(4)+in_buf[761]*(2)+in_buf[762]*(0)+in_buf[763]*(-2)+in_buf[764]*(5)+in_buf[765]*(21)+in_buf[766]*(24)+in_buf[767]*(45)+in_buf[768]*(14)+in_buf[769]*(17)+in_buf[770]*(23)+in_buf[771]*(16)+in_buf[772]*(9)+in_buf[773]*(5)+in_buf[774]*(0)+in_buf[775]*(-1)+in_buf[776]*(1)+in_buf[777]*(-23)+in_buf[778]*(-29)+in_buf[779]*(4)+in_buf[780]*(-2)+in_buf[781]*(2)+in_buf[782]*(-3)+in_buf[783]*(4);
assign in_buf_weight027=in_buf[0]*(3)+in_buf[1]*(-3)+in_buf[2]*(5)+in_buf[3]*(-1)+in_buf[4]*(-2)+in_buf[5]*(-1)+in_buf[6]*(2)+in_buf[7]*(4)+in_buf[8]*(-1)+in_buf[9]*(-3)+in_buf[10]*(0)+in_buf[11]*(4)+in_buf[12]*(-1)+in_buf[13]*(-3)+in_buf[14]*(3)+in_buf[15]*(0)+in_buf[16]*(0)+in_buf[17]*(2)+in_buf[18]*(-3)+in_buf[19]*(-3)+in_buf[20]*(2)+in_buf[21]*(0)+in_buf[22]*(-2)+in_buf[23]*(2)+in_buf[24]*(0)+in_buf[25]*(4)+in_buf[26]*(-1)+in_buf[27]*(0)+in_buf[28]*(3)+in_buf[29]*(0)+in_buf[30]*(2)+in_buf[31]*(-1)+in_buf[32]*(3)+in_buf[33]*(0)+in_buf[34]*(0)+in_buf[35]*(3)+in_buf[36]*(1)+in_buf[37]*(0)+in_buf[38]*(-1)+in_buf[39]*(-1)+in_buf[40]*(2)+in_buf[41]*(2)+in_buf[42]*(-3)+in_buf[43]*(1)+in_buf[44]*(-2)+in_buf[45]*(1)+in_buf[46]*(2)+in_buf[47]*(-1)+in_buf[48]*(0)+in_buf[49]*(-3)+in_buf[50]*(2)+in_buf[51]*(1)+in_buf[52]*(1)+in_buf[53]*(2)+in_buf[54]*(2)+in_buf[55]*(0)+in_buf[56]*(0)+in_buf[57]*(3)+in_buf[58]*(2)+in_buf[59]*(-1)+in_buf[60]*(-3)+in_buf[61]*(1)+in_buf[62]*(-2)+in_buf[63]*(0)+in_buf[64]*(3)+in_buf[65]*(-1)+in_buf[66]*(0)+in_buf[67]*(2)+in_buf[68]*(1)+in_buf[69]*(-4)+in_buf[70]*(-2)+in_buf[71]*(-2)+in_buf[72]*(1)+in_buf[73]*(3)+in_buf[74]*(2)+in_buf[75]*(-3)+in_buf[76]*(-1)+in_buf[77]*(-1)+in_buf[78]*(-2)+in_buf[79]*(0)+in_buf[80]*(4)+in_buf[81]*(3)+in_buf[82]*(-1)+in_buf[83]*(0)+in_buf[84]*(0)+in_buf[85]*(-4)+in_buf[86]*(-3)+in_buf[87]*(5)+in_buf[88]*(0)+in_buf[89]*(3)+in_buf[90]*(3)+in_buf[91]*(3)+in_buf[92]*(-1)+in_buf[93]*(0)+in_buf[94]*(0)+in_buf[95]*(1)+in_buf[96]*(-1)+in_buf[97]*(2)+in_buf[98]*(2)+in_buf[99]*(1)+in_buf[100]*(3)+in_buf[101]*(0)+in_buf[102]*(2)+in_buf[103]*(3)+in_buf[104]*(2)+in_buf[105]*(3)+in_buf[106]*(0)+in_buf[107]*(0)+in_buf[108]*(0)+in_buf[109]*(1)+in_buf[110]*(-1)+in_buf[111]*(-1)+in_buf[112]*(-2)+in_buf[113]*(-3)+in_buf[114]*(4)+in_buf[115]*(3)+in_buf[116]*(3)+in_buf[117]*(0)+in_buf[118]*(2)+in_buf[119]*(1)+in_buf[120]*(4)+in_buf[121]*(0)+in_buf[122]*(0)+in_buf[123]*(2)+in_buf[124]*(2)+in_buf[125]*(3)+in_buf[126]*(3)+in_buf[127]*(0)+in_buf[128]*(0)+in_buf[129]*(-1)+in_buf[130]*(1)+in_buf[131]*(4)+in_buf[132]*(4)+in_buf[133]*(0)+in_buf[134]*(0)+in_buf[135]*(2)+in_buf[136]*(-3)+in_buf[137]*(0)+in_buf[138]*(2)+in_buf[139]*(-2)+in_buf[140]*(0)+in_buf[141]*(0)+in_buf[142]*(-2)+in_buf[143]*(3)+in_buf[144]*(2)+in_buf[145]*(0)+in_buf[146]*(-1)+in_buf[147]*(2)+in_buf[148]*(0)+in_buf[149]*(-1)+in_buf[150]*(0)+in_buf[151]*(3)+in_buf[152]*(0)+in_buf[153]*(0)+in_buf[154]*(2)+in_buf[155]*(0)+in_buf[156]*(-3)+in_buf[157]*(-2)+in_buf[158]*(3)+in_buf[159]*(-1)+in_buf[160]*(-2)+in_buf[161]*(-1)+in_buf[162]*(0)+in_buf[163]*(-3)+in_buf[164]*(1)+in_buf[165]*(2)+in_buf[166]*(4)+in_buf[167]*(-1)+in_buf[168]*(3)+in_buf[169]*(-1)+in_buf[170]*(0)+in_buf[171]*(3)+in_buf[172]*(2)+in_buf[173]*(2)+in_buf[174]*(3)+in_buf[175]*(0)+in_buf[176]*(2)+in_buf[177]*(0)+in_buf[178]*(-2)+in_buf[179]*(3)+in_buf[180]*(-5)+in_buf[181]*(1)+in_buf[182]*(0)+in_buf[183]*(3)+in_buf[184]*(-4)+in_buf[185]*(-3)+in_buf[186]*(3)+in_buf[187]*(0)+in_buf[188]*(-1)+in_buf[189]*(1)+in_buf[190]*(1)+in_buf[191]*(-3)+in_buf[192]*(4)+in_buf[193]*(0)+in_buf[194]*(0)+in_buf[195]*(3)+in_buf[196]*(0)+in_buf[197]*(-1)+in_buf[198]*(4)+in_buf[199]*(3)+in_buf[200]*(1)+in_buf[201]*(0)+in_buf[202]*(0)+in_buf[203]*(-3)+in_buf[204]*(0)+in_buf[205]*(-4)+in_buf[206]*(-3)+in_buf[207]*(-3)+in_buf[208]*(-3)+in_buf[209]*(0)+in_buf[210]*(-1)+in_buf[211]*(1)+in_buf[212]*(2)+in_buf[213]*(-4)+in_buf[214]*(-1)+in_buf[215]*(2)+in_buf[216]*(2)+in_buf[217]*(0)+in_buf[218]*(0)+in_buf[219]*(0)+in_buf[220]*(-3)+in_buf[221]*(1)+in_buf[222]*(0)+in_buf[223]*(-3)+in_buf[224]*(4)+in_buf[225]*(2)+in_buf[226]*(3)+in_buf[227]*(1)+in_buf[228]*(3)+in_buf[229]*(-1)+in_buf[230]*(0)+in_buf[231]*(-3)+in_buf[232]*(-3)+in_buf[233]*(-2)+in_buf[234]*(-4)+in_buf[235]*(-1)+in_buf[236]*(-4)+in_buf[237]*(-3)+in_buf[238]*(-1)+in_buf[239]*(-3)+in_buf[240]*(-1)+in_buf[241]*(3)+in_buf[242]*(2)+in_buf[243]*(-3)+in_buf[244]*(1)+in_buf[245]*(0)+in_buf[246]*(-2)+in_buf[247]*(-3)+in_buf[248]*(-2)+in_buf[249]*(2)+in_buf[250]*(-3)+in_buf[251]*(4)+in_buf[252]*(-2)+in_buf[253]*(-3)+in_buf[254]*(1)+in_buf[255]*(3)+in_buf[256]*(-2)+in_buf[257]*(3)+in_buf[258]*(3)+in_buf[259]*(3)+in_buf[260]*(-2)+in_buf[261]*(-4)+in_buf[262]*(-4)+in_buf[263]*(3)+in_buf[264]*(-1)+in_buf[265]*(-1)+in_buf[266]*(0)+in_buf[267]*(-2)+in_buf[268]*(-1)+in_buf[269]*(-1)+in_buf[270]*(2)+in_buf[271]*(-4)+in_buf[272]*(1)+in_buf[273]*(0)+in_buf[274]*(1)+in_buf[275]*(-3)+in_buf[276]*(-1)+in_buf[277]*(1)+in_buf[278]*(2)+in_buf[279]*(0)+in_buf[280]*(0)+in_buf[281]*(3)+in_buf[282]*(2)+in_buf[283]*(3)+in_buf[284]*(4)+in_buf[285]*(0)+in_buf[286]*(4)+in_buf[287]*(0)+in_buf[288]*(5)+in_buf[289]*(1)+in_buf[290]*(-2)+in_buf[291]*(1)+in_buf[292]*(-1)+in_buf[293]*(-4)+in_buf[294]*(-3)+in_buf[295]*(-1)+in_buf[296]*(-4)+in_buf[297]*(-2)+in_buf[298]*(3)+in_buf[299]*(3)+in_buf[300]*(-2)+in_buf[301]*(1)+in_buf[302]*(3)+in_buf[303]*(0)+in_buf[304]*(-1)+in_buf[305]*(-3)+in_buf[306]*(-2)+in_buf[307]*(0)+in_buf[308]*(0)+in_buf[309]*(3)+in_buf[310]*(1)+in_buf[311]*(5)+in_buf[312]*(-1)+in_buf[313]*(0)+in_buf[314]*(4)+in_buf[315]*(-1)+in_buf[316]*(-1)+in_buf[317]*(-2)+in_buf[318]*(-3)+in_buf[319]*(-1)+in_buf[320]*(0)+in_buf[321]*(-3)+in_buf[322]*(-3)+in_buf[323]*(0)+in_buf[324]*(-3)+in_buf[325]*(2)+in_buf[326]*(0)+in_buf[327]*(-2)+in_buf[328]*(-1)+in_buf[329]*(-1)+in_buf[330]*(3)+in_buf[331]*(4)+in_buf[332]*(0)+in_buf[333]*(-2)+in_buf[334]*(-2)+in_buf[335]*(0)+in_buf[336]*(3)+in_buf[337]*(-1)+in_buf[338]*(-1)+in_buf[339]*(3)+in_buf[340]*(0)+in_buf[341]*(1)+in_buf[342]*(0)+in_buf[343]*(0)+in_buf[344]*(5)+in_buf[345]*(2)+in_buf[346]*(-2)+in_buf[347]*(0)+in_buf[348]*(-3)+in_buf[349]*(-1)+in_buf[350]*(-3)+in_buf[351]*(-4)+in_buf[352]*(1)+in_buf[353]*(3)+in_buf[354]*(1)+in_buf[355]*(-1)+in_buf[356]*(-4)+in_buf[357]*(0)+in_buf[358]*(0)+in_buf[359]*(-4)+in_buf[360]*(0)+in_buf[361]*(0)+in_buf[362]*(2)+in_buf[363]*(0)+in_buf[364]*(4)+in_buf[365]*(2)+in_buf[366]*(4)+in_buf[367]*(1)+in_buf[368]*(0)+in_buf[369]*(-2)+in_buf[370]*(4)+in_buf[371]*(-3)+in_buf[372]*(4)+in_buf[373]*(0)+in_buf[374]*(-1)+in_buf[375]*(0)+in_buf[376]*(-3)+in_buf[377]*(-3)+in_buf[378]*(3)+in_buf[379]*(-4)+in_buf[380]*(-2)+in_buf[381]*(-3)+in_buf[382]*(0)+in_buf[383]*(3)+in_buf[384]*(0)+in_buf[385]*(1)+in_buf[386]*(1)+in_buf[387]*(0)+in_buf[388]*(1)+in_buf[389]*(0)+in_buf[390]*(2)+in_buf[391]*(3)+in_buf[392]*(-2)+in_buf[393]*(2)+in_buf[394]*(4)+in_buf[395]*(1)+in_buf[396]*(3)+in_buf[397]*(-1)+in_buf[398]*(1)+in_buf[399]*(-2)+in_buf[400]*(-2)+in_buf[401]*(0)+in_buf[402]*(3)+in_buf[403]*(-4)+in_buf[404]*(-4)+in_buf[405]*(1)+in_buf[406]*(0)+in_buf[407]*(0)+in_buf[408]*(-3)+in_buf[409]*(0)+in_buf[410]*(-3)+in_buf[411]*(2)+in_buf[412]*(2)+in_buf[413]*(1)+in_buf[414]*(2)+in_buf[415]*(-4)+in_buf[416]*(-4)+in_buf[417]*(-2)+in_buf[418]*(2)+in_buf[419]*(-1)+in_buf[420]*(-2)+in_buf[421]*(3)+in_buf[422]*(2)+in_buf[423]*(0)+in_buf[424]*(4)+in_buf[425]*(0)+in_buf[426]*(2)+in_buf[427]*(-1)+in_buf[428]*(4)+in_buf[429]*(0)+in_buf[430]*(0)+in_buf[431]*(0)+in_buf[432]*(1)+in_buf[433]*(-2)+in_buf[434]*(0)+in_buf[435]*(-2)+in_buf[436]*(2)+in_buf[437]*(-1)+in_buf[438]*(2)+in_buf[439]*(1)+in_buf[440]*(-3)+in_buf[441]*(-5)+in_buf[442]*(-2)+in_buf[443]*(1)+in_buf[444]*(-3)+in_buf[445]*(0)+in_buf[446]*(4)+in_buf[447]*(0)+in_buf[448]*(-2)+in_buf[449]*(0)+in_buf[450]*(-1)+in_buf[451]*(1)+in_buf[452]*(5)+in_buf[453]*(-1)+in_buf[454]*(2)+in_buf[455]*(0)+in_buf[456]*(0)+in_buf[457]*(1)+in_buf[458]*(3)+in_buf[459]*(2)+in_buf[460]*(-2)+in_buf[461]*(-1)+in_buf[462]*(-1)+in_buf[463]*(-3)+in_buf[464]*(-3)+in_buf[465]*(-2)+in_buf[466]*(0)+in_buf[467]*(3)+in_buf[468]*(-2)+in_buf[469]*(2)+in_buf[470]*(-3)+in_buf[471]*(-3)+in_buf[472]*(3)+in_buf[473]*(-2)+in_buf[474]*(4)+in_buf[475]*(4)+in_buf[476]*(3)+in_buf[477]*(3)+in_buf[478]*(-2)+in_buf[479]*(-2)+in_buf[480]*(3)+in_buf[481]*(0)+in_buf[482]*(2)+in_buf[483]*(-2)+in_buf[484]*(3)+in_buf[485]*(-1)+in_buf[486]*(3)+in_buf[487]*(-2)+in_buf[488]*(-1)+in_buf[489]*(1)+in_buf[490]*(-2)+in_buf[491]*(0)+in_buf[492]*(0)+in_buf[493]*(1)+in_buf[494]*(-2)+in_buf[495]*(3)+in_buf[496]*(0)+in_buf[497]*(-2)+in_buf[498]*(0)+in_buf[499]*(-3)+in_buf[500]*(1)+in_buf[501]*(-3)+in_buf[502]*(-1)+in_buf[503]*(3)+in_buf[504]*(0)+in_buf[505]*(0)+in_buf[506]*(-2)+in_buf[507]*(1)+in_buf[508]*(-2)+in_buf[509]*(1)+in_buf[510]*(-1)+in_buf[511]*(-3)+in_buf[512]*(1)+in_buf[513]*(3)+in_buf[514]*(0)+in_buf[515]*(3)+in_buf[516]*(-2)+in_buf[517]*(0)+in_buf[518]*(-4)+in_buf[519]*(-3)+in_buf[520]*(0)+in_buf[521]*(0)+in_buf[522]*(2)+in_buf[523]*(-1)+in_buf[524]*(0)+in_buf[525]*(0)+in_buf[526]*(-3)+in_buf[527]*(3)+in_buf[528]*(-3)+in_buf[529]*(-1)+in_buf[530]*(4)+in_buf[531]*(4)+in_buf[532]*(4)+in_buf[533]*(1)+in_buf[534]*(2)+in_buf[535]*(0)+in_buf[536]*(-3)+in_buf[537]*(0)+in_buf[538]*(2)+in_buf[539]*(2)+in_buf[540]*(2)+in_buf[541]*(1)+in_buf[542]*(0)+in_buf[543]*(2)+in_buf[544]*(-2)+in_buf[545]*(3)+in_buf[546]*(-1)+in_buf[547]*(-1)+in_buf[548]*(0)+in_buf[549]*(-1)+in_buf[550]*(-2)+in_buf[551]*(-4)+in_buf[552]*(1)+in_buf[553]*(0)+in_buf[554]*(2)+in_buf[555]*(-3)+in_buf[556]*(1)+in_buf[557]*(0)+in_buf[558]*(-2)+in_buf[559]*(-2)+in_buf[560]*(4)+in_buf[561]*(2)+in_buf[562]*(0)+in_buf[563]*(3)+in_buf[564]*(0)+in_buf[565]*(-1)+in_buf[566]*(1)+in_buf[567]*(3)+in_buf[568]*(0)+in_buf[569]*(2)+in_buf[570]*(-2)+in_buf[571]*(-1)+in_buf[572]*(-1)+in_buf[573]*(-5)+in_buf[574]*(-4)+in_buf[575]*(1)+in_buf[576]*(-3)+in_buf[577]*(-1)+in_buf[578]*(0)+in_buf[579]*(3)+in_buf[580]*(-3)+in_buf[581]*(-3)+in_buf[582]*(0)+in_buf[583]*(-1)+in_buf[584]*(2)+in_buf[585]*(-1)+in_buf[586]*(0)+in_buf[587]*(-1)+in_buf[588]*(2)+in_buf[589]*(3)+in_buf[590]*(0)+in_buf[591]*(0)+in_buf[592]*(-3)+in_buf[593]*(3)+in_buf[594]*(-4)+in_buf[595]*(-4)+in_buf[596]*(1)+in_buf[597]*(3)+in_buf[598]*(-1)+in_buf[599]*(-3)+in_buf[600]*(2)+in_buf[601]*(-4)+in_buf[602]*(0)+in_buf[603]*(-4)+in_buf[604]*(0)+in_buf[605]*(0)+in_buf[606]*(0)+in_buf[607]*(-2)+in_buf[608]*(-2)+in_buf[609]*(1)+in_buf[610]*(0)+in_buf[611]*(-2)+in_buf[612]*(0)+in_buf[613]*(0)+in_buf[614]*(-1)+in_buf[615]*(1)+in_buf[616]*(-3)+in_buf[617]*(0)+in_buf[618]*(-2)+in_buf[619]*(1)+in_buf[620]*(-2)+in_buf[621]*(0)+in_buf[622]*(-1)+in_buf[623]*(-3)+in_buf[624]*(-1)+in_buf[625]*(-4)+in_buf[626]*(-4)+in_buf[627]*(2)+in_buf[628]*(-2)+in_buf[629]*(3)+in_buf[630]*(0)+in_buf[631]*(-1)+in_buf[632]*(-4)+in_buf[633]*(0)+in_buf[634]*(4)+in_buf[635]*(1)+in_buf[636]*(-1)+in_buf[637]*(0)+in_buf[638]*(-3)+in_buf[639]*(0)+in_buf[640]*(1)+in_buf[641]*(-1)+in_buf[642]*(2)+in_buf[643]*(-3)+in_buf[644]*(0)+in_buf[645]*(1)+in_buf[646]*(-1)+in_buf[647]*(4)+in_buf[648]*(3)+in_buf[649]*(2)+in_buf[650]*(-1)+in_buf[651]*(0)+in_buf[652]*(1)+in_buf[653]*(3)+in_buf[654]*(-3)+in_buf[655]*(0)+in_buf[656]*(0)+in_buf[657]*(-3)+in_buf[658]*(-2)+in_buf[659]*(-1)+in_buf[660]*(1)+in_buf[661]*(-1)+in_buf[662]*(4)+in_buf[663]*(4)+in_buf[664]*(2)+in_buf[665]*(1)+in_buf[666]*(2)+in_buf[667]*(3)+in_buf[668]*(-3)+in_buf[669]*(-2)+in_buf[670]*(-2)+in_buf[671]*(2)+in_buf[672]*(-2)+in_buf[673]*(-1)+in_buf[674]*(2)+in_buf[675]*(1)+in_buf[676]*(0)+in_buf[677]*(2)+in_buf[678]*(0)+in_buf[679]*(1)+in_buf[680]*(3)+in_buf[681]*(-1)+in_buf[682]*(-2)+in_buf[683]*(-2)+in_buf[684]*(0)+in_buf[685]*(2)+in_buf[686]*(0)+in_buf[687]*(2)+in_buf[688]*(5)+in_buf[689]*(-1)+in_buf[690]*(4)+in_buf[691]*(0)+in_buf[692]*(-3)+in_buf[693]*(5)+in_buf[694]*(4)+in_buf[695]*(0)+in_buf[696]*(1)+in_buf[697]*(-1)+in_buf[698]*(3)+in_buf[699]*(2)+in_buf[700]*(4)+in_buf[701]*(-3)+in_buf[702]*(3)+in_buf[703]*(-1)+in_buf[704]*(-3)+in_buf[705]*(4)+in_buf[706]*(3)+in_buf[707]*(1)+in_buf[708]*(2)+in_buf[709]*(1)+in_buf[710]*(-3)+in_buf[711]*(0)+in_buf[712]*(-3)+in_buf[713]*(-1)+in_buf[714]*(2)+in_buf[715]*(5)+in_buf[716]*(2)+in_buf[717]*(2)+in_buf[718]*(-2)+in_buf[719]*(4)+in_buf[720]*(0)+in_buf[721]*(0)+in_buf[722]*(-4)+in_buf[723]*(-1)+in_buf[724]*(0)+in_buf[725]*(-1)+in_buf[726]*(-1)+in_buf[727]*(2)+in_buf[728]*(1)+in_buf[729]*(0)+in_buf[730]*(0)+in_buf[731]*(-1)+in_buf[732]*(4)+in_buf[733]*(-2)+in_buf[734]*(1)+in_buf[735]*(-2)+in_buf[736]*(2)+in_buf[737]*(4)+in_buf[738]*(-3)+in_buf[739]*(0)+in_buf[740]*(4)+in_buf[741]*(1)+in_buf[742]*(-2)+in_buf[743]*(2)+in_buf[744]*(0)+in_buf[745]*(0)+in_buf[746]*(4)+in_buf[747]*(4)+in_buf[748]*(1)+in_buf[749]*(4)+in_buf[750]*(-2)+in_buf[751]*(-1)+in_buf[752]*(-2)+in_buf[753]*(0)+in_buf[754]*(-1)+in_buf[755]*(0)+in_buf[756]*(3)+in_buf[757]*(5)+in_buf[758]*(4)+in_buf[759]*(-3)+in_buf[760]*(-2)+in_buf[761]*(3)+in_buf[762]*(-3)+in_buf[763]*(-3)+in_buf[764]*(-3)+in_buf[765]*(2)+in_buf[766]*(0)+in_buf[767]*(1)+in_buf[768]*(4)+in_buf[769]*(1)+in_buf[770]*(-3)+in_buf[771]*(-1)+in_buf[772]*(2)+in_buf[773]*(2)+in_buf[774]*(0)+in_buf[775]*(1)+in_buf[776]*(0)+in_buf[777]*(4)+in_buf[778]*(-1)+in_buf[779]*(1)+in_buf[780]*(-2)+in_buf[781]*(-1)+in_buf[782]*(0)+in_buf[783]*(4);
assign in_buf_weight028=in_buf[0]*(-2)+in_buf[1]*(4)+in_buf[2]*(-2)+in_buf[3]*(4)+in_buf[4]*(-1)+in_buf[5]*(-3)+in_buf[6]*(0)+in_buf[7]*(0)+in_buf[8]*(-3)+in_buf[9]*(-1)+in_buf[10]*(1)+in_buf[11]*(2)+in_buf[12]*(11)+in_buf[13]*(9)+in_buf[14]*(0)+in_buf[15]*(1)+in_buf[16]*(4)+in_buf[17]*(3)+in_buf[18]*(2)+in_buf[19]*(0)+in_buf[20]*(2)+in_buf[21]*(0)+in_buf[22]*(2)+in_buf[23]*(2)+in_buf[24]*(0)+in_buf[25]*(4)+in_buf[26]*(-2)+in_buf[27]*(4)+in_buf[28]*(-2)+in_buf[29]*(0)+in_buf[30]*(0)+in_buf[31]*(-3)+in_buf[32]*(1)+in_buf[33]*(2)+in_buf[34]*(-2)+in_buf[35]*(-3)+in_buf[36]*(-1)+in_buf[37]*(-4)+in_buf[38]*(9)+in_buf[39]*(-11)+in_buf[40]*(-22)+in_buf[41]*(-11)+in_buf[42]*(0)+in_buf[43]*(-22)+in_buf[44]*(-40)+in_buf[45]*(-28)+in_buf[46]*(4)+in_buf[47]*(6)+in_buf[48]*(9)+in_buf[49]*(12)+in_buf[50]*(5)+in_buf[51]*(-2)+in_buf[52]*(0)+in_buf[53]*(1)+in_buf[54]*(-2)+in_buf[55]*(-1)+in_buf[56]*(0)+in_buf[57]*(0)+in_buf[58]*(-3)+in_buf[59]*(-24)+in_buf[60]*(-26)+in_buf[61]*(4)+in_buf[62]*(-4)+in_buf[63]*(-20)+in_buf[64]*(-6)+in_buf[65]*(-6)+in_buf[66]*(-21)+in_buf[67]*(-15)+in_buf[68]*(16)+in_buf[69]*(27)+in_buf[70]*(26)+in_buf[71]*(9)+in_buf[72]*(-14)+in_buf[73]*(-1)+in_buf[74]*(-3)+in_buf[75]*(7)+in_buf[76]*(11)+in_buf[77]*(1)+in_buf[78]*(1)+in_buf[79]*(4)+in_buf[80]*(-7)+in_buf[81]*(-7)+in_buf[82]*(3)+in_buf[83]*(1)+in_buf[84]*(-3)+in_buf[85]*(2)+in_buf[86]*(12)+in_buf[87]*(-32)+in_buf[88]*(-21)+in_buf[89]*(4)+in_buf[90]*(-5)+in_buf[91]*(-33)+in_buf[92]*(-32)+in_buf[93]*(-34)+in_buf[94]*(-21)+in_buf[95]*(0)+in_buf[96]*(11)+in_buf[97]*(0)+in_buf[98]*(-28)+in_buf[99]*(-44)+in_buf[100]*(-41)+in_buf[101]*(-8)+in_buf[102]*(10)+in_buf[103]*(13)+in_buf[104]*(3)+in_buf[105]*(13)+in_buf[106]*(30)+in_buf[107]*(-13)+in_buf[108]*(-32)+in_buf[109]*(16)+in_buf[110]*(14)+in_buf[111]*(-2)+in_buf[112]*(1)+in_buf[113]*(-1)+in_buf[114]*(18)+in_buf[115]*(-9)+in_buf[116]*(-28)+in_buf[117]*(-14)+in_buf[118]*(-13)+in_buf[119]*(-38)+in_buf[120]*(-32)+in_buf[121]*(-30)+in_buf[122]*(-22)+in_buf[123]*(-13)+in_buf[124]*(-18)+in_buf[125]*(-30)+in_buf[126]*(-36)+in_buf[127]*(-33)+in_buf[128]*(-23)+in_buf[129]*(-17)+in_buf[130]*(1)+in_buf[131]*(13)+in_buf[132]*(-3)+in_buf[133]*(-5)+in_buf[134]*(-4)+in_buf[135]*(47)+in_buf[136]*(27)+in_buf[137]*(19)+in_buf[138]*(6)+in_buf[139]*(3)+in_buf[140]*(-2)+in_buf[141]*(-3)+in_buf[142]*(4)+in_buf[143]*(-9)+in_buf[144]*(-10)+in_buf[145]*(-12)+in_buf[146]*(-34)+in_buf[147]*(-54)+in_buf[148]*(-30)+in_buf[149]*(-49)+in_buf[150]*(-42)+in_buf[151]*(-15)+in_buf[152]*(-7)+in_buf[153]*(-13)+in_buf[154]*(-17)+in_buf[155]*(-26)+in_buf[156]*(-38)+in_buf[157]*(-36)+in_buf[158]*(-33)+in_buf[159]*(-16)+in_buf[160]*(7)+in_buf[161]*(-3)+in_buf[162]*(-1)+in_buf[163]*(14)+in_buf[164]*(25)+in_buf[165]*(35)+in_buf[166]*(6)+in_buf[167]*(20)+in_buf[168]*(0)+in_buf[169]*(-14)+in_buf[170]*(3)+in_buf[171]*(-14)+in_buf[172]*(-11)+in_buf[173]*(-6)+in_buf[174]*(-21)+in_buf[175]*(-31)+in_buf[176]*(-51)+in_buf[177]*(-41)+in_buf[178]*(-23)+in_buf[179]*(6)+in_buf[180]*(10)+in_buf[181]*(-3)+in_buf[182]*(-6)+in_buf[183]*(-17)+in_buf[184]*(-27)+in_buf[185]*(-15)+in_buf[186]*(-2)+in_buf[187]*(7)+in_buf[188]*(11)+in_buf[189]*(15)+in_buf[190]*(27)+in_buf[191]*(18)+in_buf[192]*(40)+in_buf[193]*(55)+in_buf[194]*(17)+in_buf[195]*(-11)+in_buf[196]*(0)+in_buf[197]*(-15)+in_buf[198]*(-19)+in_buf[199]*(-11)+in_buf[200]*(-15)+in_buf[201]*(-2)+in_buf[202]*(-20)+in_buf[203]*(-34)+in_buf[204]*(-44)+in_buf[205]*(0)+in_buf[206]*(21)+in_buf[207]*(14)+in_buf[208]*(5)+in_buf[209]*(7)+in_buf[210]*(0)+in_buf[211]*(4)+in_buf[212]*(-14)+in_buf[213]*(-9)+in_buf[214]*(3)+in_buf[215]*(11)+in_buf[216]*(13)+in_buf[217]*(23)+in_buf[218]*(25)+in_buf[219]*(19)+in_buf[220]*(19)+in_buf[221]*(10)+in_buf[222]*(32)+in_buf[223]*(4)+in_buf[224]*(-30)+in_buf[225]*(-17)+in_buf[226]*(-9)+in_buf[227]*(-13)+in_buf[228]*(8)+in_buf[229]*(0)+in_buf[230]*(6)+in_buf[231]*(-3)+in_buf[232]*(0)+in_buf[233]*(11)+in_buf[234]*(12)+in_buf[235]*(4)+in_buf[236]*(1)+in_buf[237]*(1)+in_buf[238]*(-4)+in_buf[239]*(0)+in_buf[240]*(-13)+in_buf[241]*(3)+in_buf[242]*(14)+in_buf[243]*(15)+in_buf[244]*(5)+in_buf[245]*(10)+in_buf[246]*(2)+in_buf[247]*(15)+in_buf[248]*(39)+in_buf[249]*(37)+in_buf[250]*(9)+in_buf[251]*(5)+in_buf[252]*(12)+in_buf[253]*(-13)+in_buf[254]*(-27)+in_buf[255]*(-36)+in_buf[256]*(-17)+in_buf[257]*(-17)+in_buf[258]*(2)+in_buf[259]*(-10)+in_buf[260]*(-5)+in_buf[261]*(7)+in_buf[262]*(4)+in_buf[263]*(3)+in_buf[264]*(-6)+in_buf[265]*(-5)+in_buf[266]*(0)+in_buf[267]*(-2)+in_buf[268]*(10)+in_buf[269]*(10)+in_buf[270]*(22)+in_buf[271]*(-5)+in_buf[272]*(0)+in_buf[273]*(13)+in_buf[274]*(9)+in_buf[275]*(5)+in_buf[276]*(49)+in_buf[277]*(66)+in_buf[278]*(34)+in_buf[279]*(11)+in_buf[280]*(19)+in_buf[281]*(-5)+in_buf[282]*(-29)+in_buf[283]*(-41)+in_buf[284]*(-29)+in_buf[285]*(-38)+in_buf[286]*(-37)+in_buf[287]*(-13)+in_buf[288]*(1)+in_buf[289]*(20)+in_buf[290]*(18)+in_buf[291]*(6)+in_buf[292]*(10)+in_buf[293]*(3)+in_buf[294]*(10)+in_buf[295]*(15)+in_buf[296]*(9)+in_buf[297]*(5)+in_buf[298]*(11)+in_buf[299]*(6)+in_buf[300]*(2)+in_buf[301]*(23)+in_buf[302]*(8)+in_buf[303]*(10)+in_buf[304]*(55)+in_buf[305]*(81)+in_buf[306]*(20)+in_buf[307]*(-7)+in_buf[308]*(7)+in_buf[309]*(-14)+in_buf[310]*(17)+in_buf[311]*(-15)+in_buf[312]*(-25)+in_buf[313]*(-26)+in_buf[314]*(-35)+in_buf[315]*(-18)+in_buf[316]*(14)+in_buf[317]*(28)+in_buf[318]*(29)+in_buf[319]*(23)+in_buf[320]*(28)+in_buf[321]*(12)+in_buf[322]*(9)+in_buf[323]*(3)+in_buf[324]*(9)+in_buf[325]*(-11)+in_buf[326]*(0)+in_buf[327]*(-5)+in_buf[328]*(-1)+in_buf[329]*(19)+in_buf[330]*(15)+in_buf[331]*(14)+in_buf[332]*(32)+in_buf[333]*(28)+in_buf[334]*(10)+in_buf[335]*(6)+in_buf[336]*(10)+in_buf[337]*(20)+in_buf[338]*(28)+in_buf[339]*(5)+in_buf[340]*(-17)+in_buf[341]*(-31)+in_buf[342]*(-35)+in_buf[343]*(2)+in_buf[344]*(24)+in_buf[345]*(25)+in_buf[346]*(27)+in_buf[347]*(29)+in_buf[348]*(18)+in_buf[349]*(21)+in_buf[350]*(-8)+in_buf[351]*(-3)+in_buf[352]*(-2)+in_buf[353]*(-13)+in_buf[354]*(-12)+in_buf[355]*(-14)+in_buf[356]*(10)+in_buf[357]*(18)+in_buf[358]*(2)+in_buf[359]*(15)+in_buf[360]*(23)+in_buf[361]*(15)+in_buf[362]*(-2)+in_buf[363]*(-17)+in_buf[364]*(13)+in_buf[365]*(4)+in_buf[366]*(21)+in_buf[367]*(2)+in_buf[368]*(-29)+in_buf[369]*(-12)+in_buf[370]*(-41)+in_buf[371]*(-4)+in_buf[372]*(14)+in_buf[373]*(42)+in_buf[374]*(38)+in_buf[375]*(22)+in_buf[376]*(8)+in_buf[377]*(-6)+in_buf[378]*(5)+in_buf[379]*(17)+in_buf[380]*(-1)+in_buf[381]*(-12)+in_buf[382]*(-27)+in_buf[383]*(-13)+in_buf[384]*(25)+in_buf[385]*(6)+in_buf[386]*(9)+in_buf[387]*(1)+in_buf[388]*(2)+in_buf[389]*(-5)+in_buf[390]*(-50)+in_buf[391]*(-12)+in_buf[392]*(22)+in_buf[393]*(6)+in_buf[394]*(24)+in_buf[395]*(10)+in_buf[396]*(8)+in_buf[397]*(20)+in_buf[398]*(-36)+in_buf[399]*(-18)+in_buf[400]*(15)+in_buf[401]*(33)+in_buf[402]*(30)+in_buf[403]*(-2)+in_buf[404]*(-18)+in_buf[405]*(-4)+in_buf[406]*(18)+in_buf[407]*(8)+in_buf[408]*(6)+in_buf[409]*(-4)+in_buf[410]*(-27)+in_buf[411]*(-8)+in_buf[412]*(-3)+in_buf[413]*(-13)+in_buf[414]*(-7)+in_buf[415]*(-9)+in_buf[416]*(-16)+in_buf[417]*(-31)+in_buf[418]*(-47)+in_buf[419]*(-14)+in_buf[420]*(23)+in_buf[421]*(4)+in_buf[422]*(1)+in_buf[423]*(30)+in_buf[424]*(18)+in_buf[425]*(1)+in_buf[426]*(-4)+in_buf[427]*(-1)+in_buf[428]*(9)+in_buf[429]*(19)+in_buf[430]*(14)+in_buf[431]*(-5)+in_buf[432]*(-17)+in_buf[433]*(-1)+in_buf[434]*(24)+in_buf[435]*(4)+in_buf[436]*(-3)+in_buf[437]*(10)+in_buf[438]*(-8)+in_buf[439]*(-24)+in_buf[440]*(-17)+in_buf[441]*(-14)+in_buf[442]*(-4)+in_buf[443]*(-2)+in_buf[444]*(-25)+in_buf[445]*(-42)+in_buf[446]*(-17)+in_buf[447]*(-15)+in_buf[448]*(3)+in_buf[449]*(0)+in_buf[450]*(-15)+in_buf[451]*(34)+in_buf[452]*(2)+in_buf[453]*(-8)+in_buf[454]*(-1)+in_buf[455]*(-5)+in_buf[456]*(-10)+in_buf[457]*(0)+in_buf[458]*(-14)+in_buf[459]*(-20)+in_buf[460]*(-4)+in_buf[461]*(12)+in_buf[462]*(3)+in_buf[463]*(3)+in_buf[464]*(3)+in_buf[465]*(-6)+in_buf[466]*(-30)+in_buf[467]*(-21)+in_buf[468]*(-14)+in_buf[469]*(-4)+in_buf[470]*(-6)+in_buf[471]*(-19)+in_buf[472]*(-43)+in_buf[473]*(-49)+in_buf[474]*(-55)+in_buf[475]*(-6)+in_buf[476]*(4)+in_buf[477]*(-1)+in_buf[478]*(-21)+in_buf[479]*(-3)+in_buf[480]*(-4)+in_buf[481]*(-12)+in_buf[482]*(-5)+in_buf[483]*(-18)+in_buf[484]*(-14)+in_buf[485]*(0)+in_buf[486]*(8)+in_buf[487]*(-2)+in_buf[488]*(-4)+in_buf[489]*(10)+in_buf[490]*(14)+in_buf[491]*(10)+in_buf[492]*(4)+in_buf[493]*(-5)+in_buf[494]*(-12)+in_buf[495]*(-24)+in_buf[496]*(-2)+in_buf[497]*(-24)+in_buf[498]*(-23)+in_buf[499]*(-26)+in_buf[500]*(-34)+in_buf[501]*(-42)+in_buf[502]*(-33)+in_buf[503]*(-28)+in_buf[504]*(-15)+in_buf[505]*(0)+in_buf[506]*(-10)+in_buf[507]*(-19)+in_buf[508]*(-17)+in_buf[509]*(-30)+in_buf[510]*(-25)+in_buf[511]*(-22)+in_buf[512]*(-25)+in_buf[513]*(-4)+in_buf[514]*(-13)+in_buf[515]*(8)+in_buf[516]*(21)+in_buf[517]*(27)+in_buf[518]*(14)+in_buf[519]*(-9)+in_buf[520]*(-3)+in_buf[521]*(2)+in_buf[522]*(-10)+in_buf[523]*(-10)+in_buf[524]*(-21)+in_buf[525]*(-60)+in_buf[526]*(-52)+in_buf[527]*(-33)+in_buf[528]*(-24)+in_buf[529]*(-1)+in_buf[530]*(3)+in_buf[531]*(5)+in_buf[532]*(16)+in_buf[533]*(-6)+in_buf[534]*(-9)+in_buf[535]*(-34)+in_buf[536]*(-47)+in_buf[537]*(-66)+in_buf[538]*(-50)+in_buf[539]*(-25)+in_buf[540]*(-13)+in_buf[541]*(-10)+in_buf[542]*(-15)+in_buf[543]*(0)+in_buf[544]*(29)+in_buf[545]*(24)+in_buf[546]*(10)+in_buf[547]*(-4)+in_buf[548]*(-2)+in_buf[549]*(9)+in_buf[550]*(2)+in_buf[551]*(-16)+in_buf[552]*(-39)+in_buf[553]*(-49)+in_buf[554]*(-48)+in_buf[555]*(-50)+in_buf[556]*(-45)+in_buf[557]*(-9)+in_buf[558]*(-13)+in_buf[559]*(14)+in_buf[560]*(0)+in_buf[561]*(-2)+in_buf[562]*(-6)+in_buf[563]*(-55)+in_buf[564]*(-61)+in_buf[565]*(-50)+in_buf[566]*(-40)+in_buf[567]*(-29)+in_buf[568]*(-6)+in_buf[569]*(-5)+in_buf[570]*(4)+in_buf[571]*(5)+in_buf[572]*(28)+in_buf[573]*(7)+in_buf[574]*(1)+in_buf[575]*(-2)+in_buf[576]*(5)+in_buf[577]*(8)+in_buf[578]*(7)+in_buf[579]*(-12)+in_buf[580]*(-26)+in_buf[581]*(-37)+in_buf[582]*(-33)+in_buf[583]*(-42)+in_buf[584]*(-34)+in_buf[585]*(-12)+in_buf[586]*(-31)+in_buf[587]*(9)+in_buf[588]*(-1)+in_buf[589]*(-4)+in_buf[590]*(-16)+in_buf[591]*(-58)+in_buf[592]*(-48)+in_buf[593]*(-32)+in_buf[594]*(-23)+in_buf[595]*(-9)+in_buf[596]*(2)+in_buf[597]*(8)+in_buf[598]*(2)+in_buf[599]*(6)+in_buf[600]*(7)+in_buf[601]*(-7)+in_buf[602]*(-13)+in_buf[603]*(-5)+in_buf[604]*(-7)+in_buf[605]*(8)+in_buf[606]*(7)+in_buf[607]*(-24)+in_buf[608]*(-15)+in_buf[609]*(-16)+in_buf[610]*(-17)+in_buf[611]*(-31)+in_buf[612]*(-2)+in_buf[613]*(15)+in_buf[614]*(-32)+in_buf[615]*(-2)+in_buf[616]*(2)+in_buf[617]*(4)+in_buf[618]*(-8)+in_buf[619]*(-14)+in_buf[620]*(-35)+in_buf[621]*(-16)+in_buf[622]*(-9)+in_buf[623]*(-13)+in_buf[624]*(-10)+in_buf[625]*(4)+in_buf[626]*(16)+in_buf[627]*(8)+in_buf[628]*(0)+in_buf[629]*(3)+in_buf[630]*(4)+in_buf[631]*(-7)+in_buf[632]*(3)+in_buf[633]*(17)+in_buf[634]*(5)+in_buf[635]*(-7)+in_buf[636]*(-15)+in_buf[637]*(-10)+in_buf[638]*(-12)+in_buf[639]*(-5)+in_buf[640]*(-8)+in_buf[641]*(0)+in_buf[642]*(-17)+in_buf[643]*(-4)+in_buf[644]*(4)+in_buf[645]*(2)+in_buf[646]*(-25)+in_buf[647]*(-21)+in_buf[648]*(-24)+in_buf[649]*(-19)+in_buf[650]*(-8)+in_buf[651]*(2)+in_buf[652]*(6)+in_buf[653]*(9)+in_buf[654]*(-2)+in_buf[655]*(-4)+in_buf[656]*(18)+in_buf[657]*(4)+in_buf[658]*(6)+in_buf[659]*(-4)+in_buf[660]*(10)+in_buf[661]*(1)+in_buf[662]*(-8)+in_buf[663]*(-2)+in_buf[664]*(-22)+in_buf[665]*(-18)+in_buf[666]*(-23)+in_buf[667]*(-19)+in_buf[668]*(-28)+in_buf[669]*(-15)+in_buf[670]*(10)+in_buf[671]*(0)+in_buf[672]*(2)+in_buf[673]*(4)+in_buf[674]*(-17)+in_buf[675]*(-37)+in_buf[676]*(-59)+in_buf[677]*(-10)+in_buf[678]*(-14)+in_buf[679]*(7)+in_buf[680]*(-4)+in_buf[681]*(-3)+in_buf[682]*(-3)+in_buf[683]*(0)+in_buf[684]*(-1)+in_buf[685]*(12)+in_buf[686]*(6)+in_buf[687]*(6)+in_buf[688]*(-18)+in_buf[689]*(-31)+in_buf[690]*(-16)+in_buf[691]*(-1)+in_buf[692]*(3)+in_buf[693]*(0)+in_buf[694]*(12)+in_buf[695]*(-8)+in_buf[696]*(-9)+in_buf[697]*(7)+in_buf[698]*(-1)+in_buf[699]*(1)+in_buf[700]*(-1)+in_buf[701]*(3)+in_buf[702]*(8)+in_buf[703]*(2)+in_buf[704]*(2)+in_buf[705]*(0)+in_buf[706]*(-19)+in_buf[707]*(-20)+in_buf[708]*(-25)+in_buf[709]*(-16)+in_buf[710]*(-14)+in_buf[711]*(-4)+in_buf[712]*(-1)+in_buf[713]*(6)+in_buf[714]*(-1)+in_buf[715]*(-3)+in_buf[716]*(-26)+in_buf[717]*(-18)+in_buf[718]*(-20)+in_buf[719]*(-8)+in_buf[720]*(6)+in_buf[721]*(23)+in_buf[722]*(49)+in_buf[723]*(54)+in_buf[724]*(21)+in_buf[725]*(0)+in_buf[726]*(-2)+in_buf[727]*(-2)+in_buf[728]*(4)+in_buf[729]*(-1)+in_buf[730]*(-2)+in_buf[731]*(-5)+in_buf[732]*(0)+in_buf[733]*(4)+in_buf[734]*(1)+in_buf[735]*(-22)+in_buf[736]*(7)+in_buf[737]*(6)+in_buf[738]*(1)+in_buf[739]*(2)+in_buf[740]*(8)+in_buf[741]*(2)+in_buf[742]*(0)+in_buf[743]*(-5)+in_buf[744]*(-9)+in_buf[745]*(-4)+in_buf[746]*(-17)+in_buf[747]*(-7)+in_buf[748]*(-22)+in_buf[749]*(18)+in_buf[750]*(12)+in_buf[751]*(-8)+in_buf[752]*(10)+in_buf[753]*(5)+in_buf[754]*(3)+in_buf[755]*(0)+in_buf[756]*(1)+in_buf[757]*(1)+in_buf[758]*(4)+in_buf[759]*(2)+in_buf[760]*(-15)+in_buf[761]*(-1)+in_buf[762]*(-9)+in_buf[763]*(-14)+in_buf[764]*(-12)+in_buf[765]*(-2)+in_buf[766]*(11)+in_buf[767]*(-9)+in_buf[768]*(-10)+in_buf[769]*(0)+in_buf[770]*(-7)+in_buf[771]*(15)+in_buf[772]*(9)+in_buf[773]*(13)+in_buf[774]*(14)+in_buf[775]*(-2)+in_buf[776]*(12)+in_buf[777]*(18)+in_buf[778]*(14)+in_buf[779]*(10)+in_buf[780]*(2)+in_buf[781]*(-1)+in_buf[782]*(1)+in_buf[783]*(-3);
assign in_buf_weight029=in_buf[0]*(3)+in_buf[1]*(-2)+in_buf[2]*(1)+in_buf[3]*(1)+in_buf[4]*(-1)+in_buf[5]*(2)+in_buf[6]*(4)+in_buf[7]*(0)+in_buf[8]*(0)+in_buf[9]*(-2)+in_buf[10]*(0)+in_buf[11]*(-3)+in_buf[12]*(-11)+in_buf[13]*(-8)+in_buf[14]*(25)+in_buf[15]*(13)+in_buf[16]*(1)+in_buf[17]*(2)+in_buf[18]*(1)+in_buf[19]*(0)+in_buf[20]*(-1)+in_buf[21]*(3)+in_buf[22]*(-3)+in_buf[23]*(1)+in_buf[24]*(3)+in_buf[25]*(2)+in_buf[26]*(0)+in_buf[27]*(2)+in_buf[28]*(1)+in_buf[29]*(0)+in_buf[30]*(0)+in_buf[31]*(-2)+in_buf[32]*(-1)+in_buf[33]*(0)+in_buf[34]*(3)+in_buf[35]*(0)+in_buf[36]*(-4)+in_buf[37]*(1)+in_buf[38]*(-10)+in_buf[39]*(-6)+in_buf[40]*(-4)+in_buf[41]*(-24)+in_buf[42]*(-20)+in_buf[43]*(1)+in_buf[44]*(1)+in_buf[45]*(-7)+in_buf[46]*(-19)+in_buf[47]*(-12)+in_buf[48]*(-32)+in_buf[49]*(-19)+in_buf[50]*(-12)+in_buf[51]*(-2)+in_buf[52]*(-1)+in_buf[53]*(0)+in_buf[54]*(2)+in_buf[55]*(-3)+in_buf[56]*(1)+in_buf[57]*(1)+in_buf[58]*(-11)+in_buf[59]*(-1)+in_buf[60]*(-11)+in_buf[61]*(3)+in_buf[62]*(-1)+in_buf[63]*(-8)+in_buf[64]*(7)+in_buf[65]*(30)+in_buf[66]*(24)+in_buf[67]*(9)+in_buf[68]*(0)+in_buf[69]*(-12)+in_buf[70]*(18)+in_buf[71]*(44)+in_buf[72]*(13)+in_buf[73]*(2)+in_buf[74]*(22)+in_buf[75]*(18)+in_buf[76]*(16)+in_buf[77]*(-6)+in_buf[78]*(-20)+in_buf[79]*(8)+in_buf[80]*(13)+in_buf[81]*(10)+in_buf[82]*(1)+in_buf[83]*(1)+in_buf[84]*(0)+in_buf[85]*(3)+in_buf[86]*(-6)+in_buf[87]*(-2)+in_buf[88]*(16)+in_buf[89]*(25)+in_buf[90]*(30)+in_buf[91]*(26)+in_buf[92]*(49)+in_buf[93]*(23)+in_buf[94]*(27)+in_buf[95]*(22)+in_buf[96]*(28)+in_buf[97]*(28)+in_buf[98]*(16)+in_buf[99]*(13)+in_buf[100]*(8)+in_buf[101]*(0)+in_buf[102]*(10)+in_buf[103]*(9)+in_buf[104]*(19)+in_buf[105]*(20)+in_buf[106]*(-14)+in_buf[107]*(-26)+in_buf[108]*(9)+in_buf[109]*(19)+in_buf[110]*(-11)+in_buf[111]*(4)+in_buf[112]*(-3)+in_buf[113]*(3)+in_buf[114]*(19)+in_buf[115]*(30)+in_buf[116]*(8)+in_buf[117]*(29)+in_buf[118]*(31)+in_buf[119]*(41)+in_buf[120]*(27)+in_buf[121]*(17)+in_buf[122]*(28)+in_buf[123]*(27)+in_buf[124]*(31)+in_buf[125]*(13)+in_buf[126]*(8)+in_buf[127]*(18)+in_buf[128]*(28)+in_buf[129]*(26)+in_buf[130]*(20)+in_buf[131]*(9)+in_buf[132]*(0)+in_buf[133]*(8)+in_buf[134]*(-5)+in_buf[135]*(-2)+in_buf[136]*(20)+in_buf[137]*(34)+in_buf[138]*(28)+in_buf[139]*(-2)+in_buf[140]*(1)+in_buf[141]*(3)+in_buf[142]*(34)+in_buf[143]*(17)+in_buf[144]*(19)+in_buf[145]*(11)+in_buf[146]*(11)+in_buf[147]*(7)+in_buf[148]*(-10)+in_buf[149]*(-6)+in_buf[150]*(-13)+in_buf[151]*(5)+in_buf[152]*(10)+in_buf[153]*(-7)+in_buf[154]*(-8)+in_buf[155]*(-12)+in_buf[156]*(11)+in_buf[157]*(4)+in_buf[158]*(-8)+in_buf[159]*(-9)+in_buf[160]*(2)+in_buf[161]*(-3)+in_buf[162]*(2)+in_buf[163]*(4)+in_buf[164]*(2)+in_buf[165]*(23)+in_buf[166]*(20)+in_buf[167]*(0)+in_buf[168]*(-1)+in_buf[169]*(27)+in_buf[170]*(8)+in_buf[171]*(-20)+in_buf[172]*(-15)+in_buf[173]*(-17)+in_buf[174]*(-5)+in_buf[175]*(0)+in_buf[176]*(9)+in_buf[177]*(15)+in_buf[178]*(-9)+in_buf[179]*(0)+in_buf[180]*(5)+in_buf[181]*(-3)+in_buf[182]*(-8)+in_buf[183]*(-10)+in_buf[184]*(-1)+in_buf[185]*(5)+in_buf[186]*(2)+in_buf[187]*(5)+in_buf[188]*(6)+in_buf[189]*(-14)+in_buf[190]*(1)+in_buf[191]*(13)+in_buf[192]*(18)+in_buf[193]*(31)+in_buf[194]*(24)+in_buf[195]*(-17)+in_buf[196]*(0)+in_buf[197]*(31)+in_buf[198]*(-4)+in_buf[199]*(-27)+in_buf[200]*(-7)+in_buf[201]*(-8)+in_buf[202]*(-11)+in_buf[203]*(-7)+in_buf[204]*(22)+in_buf[205]*(3)+in_buf[206]*(9)+in_buf[207]*(7)+in_buf[208]*(11)+in_buf[209]*(7)+in_buf[210]*(-2)+in_buf[211]*(-7)+in_buf[212]*(0)+in_buf[213]*(0)+in_buf[214]*(-2)+in_buf[215]*(9)+in_buf[216]*(1)+in_buf[217]*(-8)+in_buf[218]*(-13)+in_buf[219]*(-18)+in_buf[220]*(25)+in_buf[221]*(56)+in_buf[222]*(1)+in_buf[223]*(-11)+in_buf[224]*(-13)+in_buf[225]*(0)+in_buf[226]*(3)+in_buf[227]*(13)+in_buf[228]*(-7)+in_buf[229]*(-7)+in_buf[230]*(-21)+in_buf[231]*(-7)+in_buf[232]*(-13)+in_buf[233]*(-4)+in_buf[234]*(0)+in_buf[235]*(19)+in_buf[236]*(19)+in_buf[237]*(15)+in_buf[238]*(1)+in_buf[239]*(0)+in_buf[240]*(-6)+in_buf[241]*(-11)+in_buf[242]*(-5)+in_buf[243]*(2)+in_buf[244]*(4)+in_buf[245]*(-4)+in_buf[246]*(-11)+in_buf[247]*(-6)+in_buf[248]*(22)+in_buf[249]*(37)+in_buf[250]*(6)+in_buf[251]*(28)+in_buf[252]*(-2)+in_buf[253]*(-10)+in_buf[254]*(6)+in_buf[255]*(19)+in_buf[256]*(-8)+in_buf[257]*(-15)+in_buf[258]*(-15)+in_buf[259]*(-9)+in_buf[260]*(4)+in_buf[261]*(2)+in_buf[262]*(8)+in_buf[263]*(21)+in_buf[264]*(17)+in_buf[265]*(1)+in_buf[266]*(-7)+in_buf[267]*(-22)+in_buf[268]*(-29)+in_buf[269]*(-14)+in_buf[270]*(-10)+in_buf[271]*(9)+in_buf[272]*(11)+in_buf[273]*(3)+in_buf[274]*(8)+in_buf[275]*(11)+in_buf[276]*(6)+in_buf[277]*(22)+in_buf[278]*(16)+in_buf[279]*(-16)+in_buf[280]*(-13)+in_buf[281]*(0)+in_buf[282]*(-13)+in_buf[283]*(18)+in_buf[284]*(19)+in_buf[285]*(-3)+in_buf[286]*(-1)+in_buf[287]*(12)+in_buf[288]*(8)+in_buf[289]*(-2)+in_buf[290]*(10)+in_buf[291]*(10)+in_buf[292]*(9)+in_buf[293]*(-18)+in_buf[294]*(-30)+in_buf[295]*(-50)+in_buf[296]*(-44)+in_buf[297]*(-32)+in_buf[298]*(-11)+in_buf[299]*(17)+in_buf[300]*(20)+in_buf[301]*(0)+in_buf[302]*(12)+in_buf[303]*(30)+in_buf[304]*(0)+in_buf[305]*(15)+in_buf[306]*(26)+in_buf[307]*(-5)+in_buf[308]*(-15)+in_buf[309]*(-32)+in_buf[310]*(-21)+in_buf[311]*(0)+in_buf[312]*(0)+in_buf[313]*(-5)+in_buf[314]*(-8)+in_buf[315]*(-2)+in_buf[316]*(-8)+in_buf[317]*(-6)+in_buf[318]*(-10)+in_buf[319]*(-18)+in_buf[320]*(-11)+in_buf[321]*(-24)+in_buf[322]*(-25)+in_buf[323]*(-28)+in_buf[324]*(-22)+in_buf[325]*(-10)+in_buf[326]*(-3)+in_buf[327]*(20)+in_buf[328]*(12)+in_buf[329]*(-10)+in_buf[330]*(-8)+in_buf[331]*(-2)+in_buf[332]*(26)+in_buf[333]*(40)+in_buf[334]*(43)+in_buf[335]*(-30)+in_buf[336]*(-22)+in_buf[337]*(-10)+in_buf[338]*(0)+in_buf[339]*(-20)+in_buf[340]*(-14)+in_buf[341]*(-16)+in_buf[342]*(-12)+in_buf[343]*(1)+in_buf[344]*(-9)+in_buf[345]*(-11)+in_buf[346]*(-2)+in_buf[347]*(-27)+in_buf[348]*(-9)+in_buf[349]*(16)+in_buf[350]*(11)+in_buf[351]*(0)+in_buf[352]*(-2)+in_buf[353]*(8)+in_buf[354]*(13)+in_buf[355]*(26)+in_buf[356]*(8)+in_buf[357]*(-3)+in_buf[358]*(-19)+in_buf[359]*(-24)+in_buf[360]*(-7)+in_buf[361]*(10)+in_buf[362]*(5)+in_buf[363]*(-21)+in_buf[364]*(9)+in_buf[365]*(-10)+in_buf[366]*(-15)+in_buf[367]*(-14)+in_buf[368]*(-35)+in_buf[369]*(-10)+in_buf[370]*(-7)+in_buf[371]*(10)+in_buf[372]*(4)+in_buf[373]*(1)+in_buf[374]*(-3)+in_buf[375]*(7)+in_buf[376]*(25)+in_buf[377]*(51)+in_buf[378]*(47)+in_buf[379]*(35)+in_buf[380]*(24)+in_buf[381]*(19)+in_buf[382]*(4)+in_buf[383]*(13)+in_buf[384]*(9)+in_buf[385]*(-7)+in_buf[386]*(-21)+in_buf[387]*(-26)+in_buf[388]*(-9)+in_buf[389]*(-2)+in_buf[390]*(48)+in_buf[391]*(27)+in_buf[392]*(21)+in_buf[393]*(-5)+in_buf[394]*(-18)+in_buf[395]*(4)+in_buf[396]*(-25)+in_buf[397]*(-8)+in_buf[398]*(8)+in_buf[399]*(-1)+in_buf[400]*(11)+in_buf[401]*(12)+in_buf[402]*(14)+in_buf[403]*(15)+in_buf[404]*(33)+in_buf[405]*(54)+in_buf[406]*(62)+in_buf[407]*(46)+in_buf[408]*(37)+in_buf[409]*(14)+in_buf[410]*(0)+in_buf[411]*(-6)+in_buf[412]*(-14)+in_buf[413]*(-16)+in_buf[414]*(-16)+in_buf[415]*(-13)+in_buf[416]*(0)+in_buf[417]*(-16)+in_buf[418]*(31)+in_buf[419]*(20)+in_buf[420]*(10)+in_buf[421]*(17)+in_buf[422]*(22)+in_buf[423]*(5)+in_buf[424]*(13)+in_buf[425]*(23)+in_buf[426]*(13)+in_buf[427]*(-2)+in_buf[428]*(0)+in_buf[429]*(4)+in_buf[430]*(11)+in_buf[431]*(19)+in_buf[432]*(31)+in_buf[433]*(57)+in_buf[434]*(44)+in_buf[435]*(36)+in_buf[436]*(27)+in_buf[437]*(4)+in_buf[438]*(1)+in_buf[439]*(-6)+in_buf[440]*(-10)+in_buf[441]*(-12)+in_buf[442]*(-9)+in_buf[443]*(1)+in_buf[444]*(12)+in_buf[445]*(-3)+in_buf[446]*(3)+in_buf[447]*(24)+in_buf[448]*(-4)+in_buf[449]*(19)+in_buf[450]*(16)+in_buf[451]*(37)+in_buf[452]*(36)+in_buf[453]*(23)+in_buf[454]*(19)+in_buf[455]*(-4)+in_buf[456]*(-11)+in_buf[457]*(0)+in_buf[458]*(3)+in_buf[459]*(9)+in_buf[460]*(25)+in_buf[461]*(35)+in_buf[462]*(32)+in_buf[463]*(15)+in_buf[464]*(14)+in_buf[465]*(6)+in_buf[466]*(0)+in_buf[467]*(0)+in_buf[468]*(-8)+in_buf[469]*(7)+in_buf[470]*(6)+in_buf[471]*(5)+in_buf[472]*(7)+in_buf[473]*(1)+in_buf[474]*(17)+in_buf[475]*(15)+in_buf[476]*(4)+in_buf[477]*(21)+in_buf[478]*(1)+in_buf[479]*(71)+in_buf[480]*(31)+in_buf[481]*(25)+in_buf[482]*(21)+in_buf[483]*(-4)+in_buf[484]*(-7)+in_buf[485]*(-12)+in_buf[486]*(-16)+in_buf[487]*(-10)+in_buf[488]*(0)+in_buf[489]*(3)+in_buf[490]*(-8)+in_buf[491]*(-2)+in_buf[492]*(9)+in_buf[493]*(4)+in_buf[494]*(-2)+in_buf[495]*(-3)+in_buf[496]*(-7)+in_buf[497]*(19)+in_buf[498]*(0)+in_buf[499]*(0)+in_buf[500]*(0)+in_buf[501]*(-23)+in_buf[502]*(23)+in_buf[503]*(19)+in_buf[504]*(-9)+in_buf[505]*(16)+in_buf[506]*(8)+in_buf[507]*(70)+in_buf[508]*(26)+in_buf[509]*(32)+in_buf[510]*(37)+in_buf[511]*(3)+in_buf[512]*(-8)+in_buf[513]*(-10)+in_buf[514]*(-3)+in_buf[515]*(-13)+in_buf[516]*(-13)+in_buf[517]*(-15)+in_buf[518]*(-10)+in_buf[519]*(1)+in_buf[520]*(7)+in_buf[521]*(2)+in_buf[522]*(-7)+in_buf[523]*(0)+in_buf[524]*(4)+in_buf[525]*(9)+in_buf[526]*(15)+in_buf[527]*(6)+in_buf[528]*(17)+in_buf[529]*(-2)+in_buf[530]*(0)+in_buf[531]*(13)+in_buf[532]*(10)+in_buf[533]*(-33)+in_buf[534]*(0)+in_buf[535]*(20)+in_buf[536]*(19)+in_buf[537]*(29)+in_buf[538]*(20)+in_buf[539]*(13)+in_buf[540]*(-3)+in_buf[541]*(-14)+in_buf[542]*(5)+in_buf[543]*(-18)+in_buf[544]*(-37)+in_buf[545]*(-12)+in_buf[546]*(-4)+in_buf[547]*(0)+in_buf[548]*(9)+in_buf[549]*(5)+in_buf[550]*(1)+in_buf[551]*(11)+in_buf[552]*(14)+in_buf[553]*(0)+in_buf[554]*(14)+in_buf[555]*(26)+in_buf[556]*(5)+in_buf[557]*(19)+in_buf[558]*(46)+in_buf[559]*(3)+in_buf[560]*(0)+in_buf[561]*(-10)+in_buf[562]*(8)+in_buf[563]*(18)+in_buf[564]*(13)+in_buf[565]*(8)+in_buf[566]*(17)+in_buf[567]*(17)+in_buf[568]*(1)+in_buf[569]*(-6)+in_buf[570]*(-1)+in_buf[571]*(-14)+in_buf[572]*(-48)+in_buf[573]*(-18)+in_buf[574]*(-5)+in_buf[575]*(0)+in_buf[576]*(4)+in_buf[577]*(5)+in_buf[578]*(12)+in_buf[579]*(11)+in_buf[580]*(16)+in_buf[581]*(10)+in_buf[582]*(12)+in_buf[583]*(16)+in_buf[584]*(-13)+in_buf[585]*(19)+in_buf[586]*(27)+in_buf[587]*(3)+in_buf[588]*(-11)+in_buf[589]*(5)+in_buf[590]*(16)+in_buf[591]*(18)+in_buf[592]*(-9)+in_buf[593]*(-20)+in_buf[594]*(0)+in_buf[595]*(5)+in_buf[596]*(0)+in_buf[597]*(-12)+in_buf[598]*(-13)+in_buf[599]*(-5)+in_buf[600]*(-19)+in_buf[601]*(-7)+in_buf[602]*(-2)+in_buf[603]*(4)+in_buf[604]*(-4)+in_buf[605]*(0)+in_buf[606]*(9)+in_buf[607]*(17)+in_buf[608]*(13)+in_buf[609]*(12)+in_buf[610]*(3)+in_buf[611]*(-5)+in_buf[612]*(-24)+in_buf[613]*(22)+in_buf[614]*(-22)+in_buf[615]*(-5)+in_buf[616]*(-8)+in_buf[617]*(15)+in_buf[618]*(28)+in_buf[619]*(34)+in_buf[620]*(2)+in_buf[621]*(-18)+in_buf[622]*(-25)+in_buf[623]*(-11)+in_buf[624]*(-27)+in_buf[625]*(-25)+in_buf[626]*(-19)+in_buf[627]*(0)+in_buf[628]*(-14)+in_buf[629]*(-7)+in_buf[630]*(0)+in_buf[631]*(-8)+in_buf[632]*(-3)+in_buf[633]*(9)+in_buf[634]*(5)+in_buf[635]*(13)+in_buf[636]*(21)+in_buf[637]*(3)+in_buf[638]*(7)+in_buf[639]*(7)+in_buf[640]*(-3)+in_buf[641]*(33)+in_buf[642]*(13)+in_buf[643]*(-2)+in_buf[644]*(0)+in_buf[645]*(2)+in_buf[646]*(41)+in_buf[647]*(53)+in_buf[648]*(38)+in_buf[649]*(1)+in_buf[650]*(-17)+in_buf[651]*(-10)+in_buf[652]*(-8)+in_buf[653]*(-14)+in_buf[654]*(-15)+in_buf[655]*(-8)+in_buf[656]*(-13)+in_buf[657]*(4)+in_buf[658]*(-7)+in_buf[659]*(-7)+in_buf[660]*(0)+in_buf[661]*(1)+in_buf[662]*(8)+in_buf[663]*(1)+in_buf[664]*(8)+in_buf[665]*(2)+in_buf[666]*(14)+in_buf[667]*(8)+in_buf[668]*(11)+in_buf[669]*(36)+in_buf[670]*(24)+in_buf[671]*(4)+in_buf[672]*(3)+in_buf[673]*(2)+in_buf[674]*(18)+in_buf[675]*(36)+in_buf[676]*(15)+in_buf[677]*(-9)+in_buf[678]*(10)+in_buf[679]*(10)+in_buf[680]*(9)+in_buf[681]*(14)+in_buf[682]*(4)+in_buf[683]*(1)+in_buf[684]*(1)+in_buf[685]*(4)+in_buf[686]*(3)+in_buf[687]*(-11)+in_buf[688]*(18)+in_buf[689]*(13)+in_buf[690]*(24)+in_buf[691]*(20)+in_buf[692]*(20)+in_buf[693]*(24)+in_buf[694]*(0)+in_buf[695]*(0)+in_buf[696]*(6)+in_buf[697]*(-13)+in_buf[698]*(-9)+in_buf[699]*(0)+in_buf[700]*(4)+in_buf[701]*(-1)+in_buf[702]*(0)+in_buf[703]*(-29)+in_buf[704]*(-14)+in_buf[705]*(9)+in_buf[706]*(33)+in_buf[707]*(46)+in_buf[708]*(44)+in_buf[709]*(45)+in_buf[710]*(51)+in_buf[711]*(25)+in_buf[712]*(48)+in_buf[713]*(54)+in_buf[714]*(32)+in_buf[715]*(28)+in_buf[716]*(44)+in_buf[717]*(56)+in_buf[718]*(45)+in_buf[719]*(41)+in_buf[720]*(26)+in_buf[721]*(14)+in_buf[722]*(14)+in_buf[723]*(29)+in_buf[724]*(40)+in_buf[725]*(-11)+in_buf[726]*(2)+in_buf[727]*(1)+in_buf[728]*(-2)+in_buf[729]*(-3)+in_buf[730]*(-1)+in_buf[731]*(-8)+in_buf[732]*(21)+in_buf[733]*(25)+in_buf[734]*(17)+in_buf[735]*(26)+in_buf[736]*(13)+in_buf[737]*(1)+in_buf[738]*(11)+in_buf[739]*(11)+in_buf[740]*(14)+in_buf[741]*(8)+in_buf[742]*(13)+in_buf[743]*(21)+in_buf[744]*(35)+in_buf[745]*(47)+in_buf[746]*(39)+in_buf[747]*(10)+in_buf[748]*(5)+in_buf[749]*(-1)+in_buf[750]*(3)+in_buf[751]*(28)+in_buf[752]*(6)+in_buf[753]*(-3)+in_buf[754]*(2)+in_buf[755]*(1)+in_buf[756]*(1)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(3)+in_buf[760]*(-17)+in_buf[761]*(-13)+in_buf[762]*(11)+in_buf[763]*(15)+in_buf[764]*(3)+in_buf[765]*(-4)+in_buf[766]*(-20)+in_buf[767]*(2)+in_buf[768]*(5)+in_buf[769]*(-12)+in_buf[770]*(17)+in_buf[771]*(25)+in_buf[772]*(-7)+in_buf[773]*(-22)+in_buf[774]*(-31)+in_buf[775]*(-22)+in_buf[776]*(-28)+in_buf[777]*(-24)+in_buf[778]*(-18)+in_buf[779]*(2)+in_buf[780]*(1)+in_buf[781]*(4)+in_buf[782]*(2)+in_buf[783]*(2);
assign in_buf_weight030=in_buf[0]*(2)+in_buf[1]*(-1)+in_buf[2]*(-2)+in_buf[3]*(2)+in_buf[4]*(0)+in_buf[5]*(4)+in_buf[6]*(4)+in_buf[7]*(1)+in_buf[8]*(3)+in_buf[9]*(3)+in_buf[10]*(4)+in_buf[11]*(-2)+in_buf[12]*(-2)+in_buf[13]*(7)+in_buf[14]*(7)+in_buf[15]*(1)+in_buf[16]*(1)+in_buf[17]*(3)+in_buf[18]*(-2)+in_buf[19]*(3)+in_buf[20]*(5)+in_buf[21]*(1)+in_buf[22]*(4)+in_buf[23]*(-1)+in_buf[24]*(3)+in_buf[25]*(0)+in_buf[26]*(-1)+in_buf[27]*(-1)+in_buf[28]*(0)+in_buf[29]*(0)+in_buf[30]*(-3)+in_buf[31]*(-2)+in_buf[32]*(3)+in_buf[33]*(0)+in_buf[34]*(-2)+in_buf[35]*(0)+in_buf[36]*(-5)+in_buf[37]*(0)+in_buf[38]*(-13)+in_buf[39]*(15)+in_buf[40]*(22)+in_buf[41]*(25)+in_buf[42]*(-10)+in_buf[43]*(12)+in_buf[44]*(27)+in_buf[45]*(24)+in_buf[46]*(0)+in_buf[47]*(-3)+in_buf[48]*(-10)+in_buf[49]*(-5)+in_buf[50]*(-7)+in_buf[51]*(-7)+in_buf[52]*(0)+in_buf[53]*(-3)+in_buf[54]*(-3)+in_buf[55]*(0)+in_buf[56]*(0)+in_buf[57]*(3)+in_buf[58]*(2)+in_buf[59]*(32)+in_buf[60]*(30)+in_buf[61]*(1)+in_buf[62]*(0)+in_buf[63]*(4)+in_buf[64]*(-18)+in_buf[65]*(-15)+in_buf[66]*(0)+in_buf[67]*(7)+in_buf[68]*(-6)+in_buf[69]*(-20)+in_buf[70]*(-18)+in_buf[71]*(-32)+in_buf[72]*(-13)+in_buf[73]*(-32)+in_buf[74]*(-31)+in_buf[75]*(-17)+in_buf[76]*(-35)+in_buf[77]*(-35)+in_buf[78]*(-18)+in_buf[79]*(-11)+in_buf[80]*(-3)+in_buf[81]*(-5)+in_buf[82]*(-1)+in_buf[83]*(3)+in_buf[84]*(-1)+in_buf[85]*(3)+in_buf[86]*(-7)+in_buf[87]*(31)+in_buf[88]*(0)+in_buf[89]*(6)+in_buf[90]*(-19)+in_buf[91]*(-3)+in_buf[92]*(-14)+in_buf[93]*(-15)+in_buf[94]*(-26)+in_buf[95]*(-3)+in_buf[96]*(8)+in_buf[97]*(-3)+in_buf[98]*(20)+in_buf[99]*(0)+in_buf[100]*(1)+in_buf[101]*(9)+in_buf[102]*(-16)+in_buf[103]*(-11)+in_buf[104]*(18)+in_buf[105]*(0)+in_buf[106]*(-26)+in_buf[107]*(-35)+in_buf[108]*(-9)+in_buf[109]*(36)+in_buf[110]*(29)+in_buf[111]*(-3)+in_buf[112]*(-1)+in_buf[113]*(7)+in_buf[114]*(2)+in_buf[115]*(11)+in_buf[116]*(35)+in_buf[117]*(12)+in_buf[118]*(-1)+in_buf[119]*(-20)+in_buf[120]*(-5)+in_buf[121]*(-6)+in_buf[122]*(-2)+in_buf[123]*(-3)+in_buf[124]*(2)+in_buf[125]*(-2)+in_buf[126]*(-2)+in_buf[127]*(6)+in_buf[128]*(6)+in_buf[129]*(12)+in_buf[130]*(10)+in_buf[131]*(8)+in_buf[132]*(6)+in_buf[133]*(-1)+in_buf[134]*(15)+in_buf[135]*(-22)+in_buf[136]*(-21)+in_buf[137]*(-9)+in_buf[138]*(-17)+in_buf[139]*(9)+in_buf[140]*(-1)+in_buf[141]*(-2)+in_buf[142]*(-10)+in_buf[143]*(1)+in_buf[144]*(31)+in_buf[145]*(30)+in_buf[146]*(3)+in_buf[147]*(-15)+in_buf[148]*(2)+in_buf[149]*(4)+in_buf[150]*(9)+in_buf[151]*(5)+in_buf[152]*(3)+in_buf[153]*(7)+in_buf[154]*(5)+in_buf[155]*(5)+in_buf[156]*(-4)+in_buf[157]*(-8)+in_buf[158]*(9)+in_buf[159]*(4)+in_buf[160]*(-3)+in_buf[161]*(-12)+in_buf[162]*(12)+in_buf[163]*(17)+in_buf[164]*(3)+in_buf[165]*(-19)+in_buf[166]*(-30)+in_buf[167]*(1)+in_buf[168]*(-3)+in_buf[169]*(27)+in_buf[170]*(23)+in_buf[171]*(38)+in_buf[172]*(39)+in_buf[173]*(22)+in_buf[174]*(8)+in_buf[175]*(6)+in_buf[176]*(21)+in_buf[177]*(17)+in_buf[178]*(20)+in_buf[179]*(11)+in_buf[180]*(12)+in_buf[181]*(21)+in_buf[182]*(3)+in_buf[183]*(-8)+in_buf[184]*(-4)+in_buf[185]*(-6)+in_buf[186]*(3)+in_buf[187]*(-2)+in_buf[188]*(0)+in_buf[189]*(17)+in_buf[190]*(9)+in_buf[191]*(11)+in_buf[192]*(9)+in_buf[193]*(-42)+in_buf[194]*(0)+in_buf[195]*(8)+in_buf[196]*(1)+in_buf[197]*(46)+in_buf[198]*(10)+in_buf[199]*(51)+in_buf[200]*(13)+in_buf[201]*(-14)+in_buf[202]*(-13)+in_buf[203]*(-1)+in_buf[204]*(14)+in_buf[205]*(9)+in_buf[206]*(1)+in_buf[207]*(-2)+in_buf[208]*(-2)+in_buf[209]*(-1)+in_buf[210]*(9)+in_buf[211]*(-1)+in_buf[212]*(8)+in_buf[213]*(5)+in_buf[214]*(3)+in_buf[215]*(-9)+in_buf[216]*(8)+in_buf[217]*(5)+in_buf[218]*(8)+in_buf[219]*(15)+in_buf[220]*(7)+in_buf[221]*(1)+in_buf[222]*(5)+in_buf[223]*(19)+in_buf[224]*(38)+in_buf[225]*(41)+in_buf[226]*(3)+in_buf[227]*(36)+in_buf[228]*(-14)+in_buf[229]*(-28)+in_buf[230]*(-18)+in_buf[231]*(-6)+in_buf[232]*(-12)+in_buf[233]*(-14)+in_buf[234]*(-23)+in_buf[235]*(-32)+in_buf[236]*(-27)+in_buf[237]*(-25)+in_buf[238]*(-3)+in_buf[239]*(6)+in_buf[240]*(12)+in_buf[241]*(2)+in_buf[242]*(1)+in_buf[243]*(-9)+in_buf[244]*(-1)+in_buf[245]*(0)+in_buf[246]*(15)+in_buf[247]*(-2)+in_buf[248]*(-16)+in_buf[249]*(-16)+in_buf[250]*(9)+in_buf[251]*(2)+in_buf[252]*(13)+in_buf[253]*(36)+in_buf[254]*(-11)+in_buf[255]*(10)+in_buf[256]*(-30)+in_buf[257]*(-28)+in_buf[258]*(-25)+in_buf[259]*(-20)+in_buf[260]*(-27)+in_buf[261]*(-43)+in_buf[262]*(-28)+in_buf[263]*(-47)+in_buf[264]*(-28)+in_buf[265]*(-21)+in_buf[266]*(0)+in_buf[267]*(0)+in_buf[268]*(6)+in_buf[269]*(2)+in_buf[270]*(5)+in_buf[271]*(5)+in_buf[272]*(8)+in_buf[273]*(8)+in_buf[274]*(10)+in_buf[275]*(-1)+in_buf[276]*(2)+in_buf[277]*(-30)+in_buf[278]*(-18)+in_buf[279]*(-30)+in_buf[280]*(20)+in_buf[281]*(25)+in_buf[282]*(29)+in_buf[283]*(3)+in_buf[284]*(-32)+in_buf[285]*(-33)+in_buf[286]*(-34)+in_buf[287]*(-36)+in_buf[288]*(-42)+in_buf[289]*(-44)+in_buf[290]*(-42)+in_buf[291]*(-35)+in_buf[292]*(-16)+in_buf[293]*(9)+in_buf[294]*(6)+in_buf[295]*(-1)+in_buf[296]*(6)+in_buf[297]*(4)+in_buf[298]*(7)+in_buf[299]*(12)+in_buf[300]*(22)+in_buf[301]*(10)+in_buf[302]*(17)+in_buf[303]*(-4)+in_buf[304]*(-4)+in_buf[305]*(-31)+in_buf[306]*(-38)+in_buf[307]*(-25)+in_buf[308]*(9)+in_buf[309]*(28)+in_buf[310]*(22)+in_buf[311]*(30)+in_buf[312]*(-6)+in_buf[313]*(-37)+in_buf[314]*(-34)+in_buf[315]*(-12)+in_buf[316]*(-18)+in_buf[317]*(-23)+in_buf[318]*(-12)+in_buf[319]*(4)+in_buf[320]*(19)+in_buf[321]*(39)+in_buf[322]*(13)+in_buf[323]*(0)+in_buf[324]*(-15)+in_buf[325]*(3)+in_buf[326]*(9)+in_buf[327]*(16)+in_buf[328]*(15)+in_buf[329]*(-1)+in_buf[330]*(11)+in_buf[331]*(0)+in_buf[332]*(-46)+in_buf[333]*(-51)+in_buf[334]*(-38)+in_buf[335]*(6)+in_buf[336]*(8)+in_buf[337]*(11)+in_buf[338]*(12)+in_buf[339]*(12)+in_buf[340]*(-10)+in_buf[341]*(-7)+in_buf[342]*(-8)+in_buf[343]*(13)+in_buf[344]*(7)+in_buf[345]*(12)+in_buf[346]*(17)+in_buf[347]*(41)+in_buf[348]*(59)+in_buf[349]*(41)+in_buf[350]*(23)+in_buf[351]*(1)+in_buf[352]*(-9)+in_buf[353]*(-4)+in_buf[354]*(6)+in_buf[355]*(-1)+in_buf[356]*(-7)+in_buf[357]*(-5)+in_buf[358]*(20)+in_buf[359]*(0)+in_buf[360]*(-34)+in_buf[361]*(-36)+in_buf[362]*(-21)+in_buf[363]*(1)+in_buf[364]*(-2)+in_buf[365]*(-3)+in_buf[366]*(41)+in_buf[367]*(37)+in_buf[368]*(31)+in_buf[369]*(31)+in_buf[370]*(35)+in_buf[371]*(29)+in_buf[372]*(24)+in_buf[373]*(6)+in_buf[374]*(32)+in_buf[375]*(28)+in_buf[376]*(35)+in_buf[377]*(14)+in_buf[378]*(-1)+in_buf[379]*(-13)+in_buf[380]*(-9)+in_buf[381]*(0)+in_buf[382]*(12)+in_buf[383]*(0)+in_buf[384]*(-11)+in_buf[385]*(6)+in_buf[386]*(0)+in_buf[387]*(10)+in_buf[388]*(5)+in_buf[389]*(-7)+in_buf[390]*(1)+in_buf[391]*(-13)+in_buf[392]*(-19)+in_buf[393]*(6)+in_buf[394]*(26)+in_buf[395]*(42)+in_buf[396]*(26)+in_buf[397]*(27)+in_buf[398]*(30)+in_buf[399]*(22)+in_buf[400]*(17)+in_buf[401]*(8)+in_buf[402]*(13)+in_buf[403]*(25)+in_buf[404]*(21)+in_buf[405]*(3)+in_buf[406]*(-13)+in_buf[407]*(-5)+in_buf[408]*(-14)+in_buf[409]*(5)+in_buf[410]*(13)+in_buf[411]*(2)+in_buf[412]*(2)+in_buf[413]*(4)+in_buf[414]*(4)+in_buf[415]*(12)+in_buf[416]*(2)+in_buf[417]*(-30)+in_buf[418]*(0)+in_buf[419]*(-6)+in_buf[420]*(-10)+in_buf[421]*(10)+in_buf[422]*(10)+in_buf[423]*(6)+in_buf[424]*(23)+in_buf[425]*(20)+in_buf[426]*(12)+in_buf[427]*(0)+in_buf[428]*(-16)+in_buf[429]*(-7)+in_buf[430]*(2)+in_buf[431]*(4)+in_buf[432]*(15)+in_buf[433]*(-6)+in_buf[434]*(-8)+in_buf[435]*(5)+in_buf[436]*(4)+in_buf[437]*(13)+in_buf[438]*(17)+in_buf[439]*(5)+in_buf[440]*(6)+in_buf[441]*(2)+in_buf[442]*(6)+in_buf[443]*(-4)+in_buf[444]*(4)+in_buf[445]*(-35)+in_buf[446]*(11)+in_buf[447]*(-2)+in_buf[448]*(0)+in_buf[449]*(14)+in_buf[450]*(20)+in_buf[451]*(-2)+in_buf[452]*(35)+in_buf[453]*(11)+in_buf[454]*(-12)+in_buf[455]*(-11)+in_buf[456]*(-17)+in_buf[457]*(-8)+in_buf[458]*(-10)+in_buf[459]*(-5)+in_buf[460]*(-1)+in_buf[461]*(-17)+in_buf[462]*(-13)+in_buf[463]*(7)+in_buf[464]*(10)+in_buf[465]*(19)+in_buf[466]*(9)+in_buf[467]*(6)+in_buf[468]*(8)+in_buf[469]*(3)+in_buf[470]*(-9)+in_buf[471]*(-22)+in_buf[472]*(-9)+in_buf[473]*(-40)+in_buf[474]*(-15)+in_buf[475]*(11)+in_buf[476]*(4)+in_buf[477]*(10)+in_buf[478]*(4)+in_buf[479]*(5)+in_buf[480]*(22)+in_buf[481]*(0)+in_buf[482]*(-18)+in_buf[483]*(-14)+in_buf[484]*(-26)+in_buf[485]*(-25)+in_buf[486]*(-17)+in_buf[487]*(-1)+in_buf[488]*(-8)+in_buf[489]*(-17)+in_buf[490]*(-21)+in_buf[491]*(1)+in_buf[492]*(12)+in_buf[493]*(17)+in_buf[494]*(7)+in_buf[495]*(1)+in_buf[496]*(-10)+in_buf[497]*(7)+in_buf[498]*(1)+in_buf[499]*(-13)+in_buf[500]*(-16)+in_buf[501]*(-31)+in_buf[502]*(12)+in_buf[503]*(14)+in_buf[504]*(28)+in_buf[505]*(8)+in_buf[506]*(25)+in_buf[507]*(5)+in_buf[508]*(0)+in_buf[509]*(-2)+in_buf[510]*(-7)+in_buf[511]*(-14)+in_buf[512]*(-5)+in_buf[513]*(-20)+in_buf[514]*(-13)+in_buf[515]*(4)+in_buf[516]*(-4)+in_buf[517]*(-10)+in_buf[518]*(-2)+in_buf[519]*(15)+in_buf[520]*(20)+in_buf[521]*(4)+in_buf[522]*(7)+in_buf[523]*(-8)+in_buf[524]*(-18)+in_buf[525]*(9)+in_buf[526]*(2)+in_buf[527]*(-38)+in_buf[528]*(-46)+in_buf[529]*(-14)+in_buf[530]*(13)+in_buf[531]*(-8)+in_buf[532]*(-15)+in_buf[533]*(46)+in_buf[534]*(21)+in_buf[535]*(7)+in_buf[536]*(2)+in_buf[537]*(12)+in_buf[538]*(8)+in_buf[539]*(-8)+in_buf[540]*(3)+in_buf[541]*(-10)+in_buf[542]*(-11)+in_buf[543]*(-2)+in_buf[544]*(14)+in_buf[545]*(6)+in_buf[546]*(14)+in_buf[547]*(8)+in_buf[548]*(-1)+in_buf[549]*(0)+in_buf[550]*(-7)+in_buf[551]*(-20)+in_buf[552]*(-13)+in_buf[553]*(-3)+in_buf[554]*(-22)+in_buf[555]*(-26)+in_buf[556]*(-36)+in_buf[557]*(-13)+in_buf[558]*(-13)+in_buf[559]*(-6)+in_buf[560]*(0)+in_buf[561]*(30)+in_buf[562]*(0)+in_buf[563]*(13)+in_buf[564]*(9)+in_buf[565]*(-6)+in_buf[566]*(-1)+in_buf[567]*(8)+in_buf[568]*(3)+in_buf[569]*(2)+in_buf[570]*(2)+in_buf[571]*(1)+in_buf[572]*(14)+in_buf[573]*(24)+in_buf[574]*(12)+in_buf[575]*(-3)+in_buf[576]*(-11)+in_buf[577]*(-5)+in_buf[578]*(-7)+in_buf[579]*(-21)+in_buf[580]*(-6)+in_buf[581]*(-17)+in_buf[582]*(-34)+in_buf[583]*(-57)+in_buf[584]*(-22)+in_buf[585]*(-6)+in_buf[586]*(18)+in_buf[587]*(-4)+in_buf[588]*(-3)+in_buf[589]*(2)+in_buf[590]*(-7)+in_buf[591]*(0)+in_buf[592]*(-22)+in_buf[593]*(-18)+in_buf[594]*(-2)+in_buf[595]*(6)+in_buf[596]*(14)+in_buf[597]*(0)+in_buf[598]*(-1)+in_buf[599]*(-5)+in_buf[600]*(0)+in_buf[601]*(2)+in_buf[602]*(-15)+in_buf[603]*(-13)+in_buf[604]*(-5)+in_buf[605]*(-15)+in_buf[606]*(-17)+in_buf[607]*(-17)+in_buf[608]*(-26)+in_buf[609]*(-21)+in_buf[610]*(-51)+in_buf[611]*(-45)+in_buf[612]*(-12)+in_buf[613]*(-20)+in_buf[614]*(34)+in_buf[615]*(6)+in_buf[616]*(4)+in_buf[617]*(21)+in_buf[618]*(1)+in_buf[619]*(-12)+in_buf[620]*(-27)+in_buf[621]*(-23)+in_buf[622]*(-2)+in_buf[623]*(15)+in_buf[624]*(13)+in_buf[625]*(2)+in_buf[626]*(4)+in_buf[627]*(-1)+in_buf[628]*(2)+in_buf[629]*(-10)+in_buf[630]*(-1)+in_buf[631]*(5)+in_buf[632]*(0)+in_buf[633]*(-14)+in_buf[634]*(-34)+in_buf[635]*(-18)+in_buf[636]*(-27)+in_buf[637]*(-15)+in_buf[638]*(-15)+in_buf[639]*(-6)+in_buf[640]*(-19)+in_buf[641]*(-19)+in_buf[642]*(31)+in_buf[643]*(3)+in_buf[644]*(-3)+in_buf[645]*(-3)+in_buf[646]*(39)+in_buf[647]*(-7)+in_buf[648]*(-27)+in_buf[649]*(-4)+in_buf[650]*(2)+in_buf[651]*(29)+in_buf[652]*(9)+in_buf[653]*(8)+in_buf[654]*(16)+in_buf[655]*(22)+in_buf[656]*(-5)+in_buf[657]*(-5)+in_buf[658]*(-2)+in_buf[659]*(-13)+in_buf[660]*(-18)+in_buf[661]*(-17)+in_buf[662]*(-17)+in_buf[663]*(-35)+in_buf[664]*(-34)+in_buf[665]*(-7)+in_buf[666]*(-4)+in_buf[667]*(-24)+in_buf[668]*(-9)+in_buf[669]*(-8)+in_buf[670]*(17)+in_buf[671]*(0)+in_buf[672]*(1)+in_buf[673]*(3)+in_buf[674]*(9)+in_buf[675]*(30)+in_buf[676]*(29)+in_buf[677]*(22)+in_buf[678]*(16)+in_buf[679]*(11)+in_buf[680]*(5)+in_buf[681]*(-7)+in_buf[682]*(-7)+in_buf[683]*(-4)+in_buf[684]*(-15)+in_buf[685]*(0)+in_buf[686]*(9)+in_buf[687]*(-18)+in_buf[688]*(-19)+in_buf[689]*(4)+in_buf[690]*(-6)+in_buf[691]*(-36)+in_buf[692]*(-46)+in_buf[693]*(-15)+in_buf[694]*(-8)+in_buf[695]*(-13)+in_buf[696]*(-8)+in_buf[697]*(-5)+in_buf[698]*(9)+in_buf[699]*(-2)+in_buf[700]*(3)+in_buf[701]*(0)+in_buf[702]*(7)+in_buf[703]*(17)+in_buf[704]*(42)+in_buf[705]*(36)+in_buf[706]*(23)+in_buf[707]*(22)+in_buf[708]*(2)+in_buf[709]*(-20)+in_buf[710]*(-3)+in_buf[711]*(4)+in_buf[712]*(-12)+in_buf[713]*(0)+in_buf[714]*(-5)+in_buf[715]*(-23)+in_buf[716]*(-16)+in_buf[717]*(-31)+in_buf[718]*(-29)+in_buf[719]*(-24)+in_buf[720]*(-51)+in_buf[721]*(-30)+in_buf[722]*(-21)+in_buf[723]*(5)+in_buf[724]*(13)+in_buf[725]*(4)+in_buf[726]*(1)+in_buf[727]*(-3)+in_buf[728]*(-2)+in_buf[729]*(0)+in_buf[730]*(0)+in_buf[731]*(11)+in_buf[732]*(-30)+in_buf[733]*(-29)+in_buf[734]*(-1)+in_buf[735]*(11)+in_buf[736]*(1)+in_buf[737]*(-7)+in_buf[738]*(9)+in_buf[739]*(18)+in_buf[740]*(14)+in_buf[741]*(28)+in_buf[742]*(-9)+in_buf[743]*(-16)+in_buf[744]*(-9)+in_buf[745]*(-20)+in_buf[746]*(-16)+in_buf[747]*(-7)+in_buf[748]*(-30)+in_buf[749]*(-27)+in_buf[750]*(-5)+in_buf[751]*(-5)+in_buf[752]*(-10)+in_buf[753]*(13)+in_buf[754]*(-1)+in_buf[755]*(-1)+in_buf[756]*(-1)+in_buf[757]*(-1)+in_buf[758]*(3)+in_buf[759]*(0)+in_buf[760]*(21)+in_buf[761]*(25)+in_buf[762]*(-7)+in_buf[763]*(-4)+in_buf[764]*(-6)+in_buf[765]*(5)+in_buf[766]*(4)+in_buf[767]*(-18)+in_buf[768]*(-11)+in_buf[769]*(5)+in_buf[770]*(-15)+in_buf[771]*(-16)+in_buf[772]*(16)+in_buf[773]*(31)+in_buf[774]*(8)+in_buf[775]*(9)+in_buf[776]*(5)+in_buf[777]*(0)+in_buf[778]*(6)+in_buf[779]*(3)+in_buf[780]*(2)+in_buf[781]*(4)+in_buf[782]*(4)+in_buf[783]*(3);
assign in_buf_weight031=in_buf[0]*(-2)+in_buf[1]*(3)+in_buf[2]*(4)+in_buf[3]*(1)+in_buf[4]*(0)+in_buf[5]*(2)+in_buf[6]*(0)+in_buf[7]*(-1)+in_buf[8]*(-2)+in_buf[9]*(3)+in_buf[10]*(2)+in_buf[11]*(0)+in_buf[12]*(0)+in_buf[13]*(-2)+in_buf[14]*(-6)+in_buf[15]*(-2)+in_buf[16]*(-2)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(0)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(3)+in_buf[23]*(4)+in_buf[24]*(4)+in_buf[25]*(-1)+in_buf[26]*(-2)+in_buf[27]*(-3)+in_buf[28]*(2)+in_buf[29]*(0)+in_buf[30]*(-3)+in_buf[31]*(-1)+in_buf[32]*(-5)+in_buf[33]*(-9)+in_buf[34]*(-13)+in_buf[35]*(-6)+in_buf[36]*(-13)+in_buf[37]*(-11)+in_buf[38]*(-10)+in_buf[39]*(-18)+in_buf[40]*(-14)+in_buf[41]*(1)+in_buf[42]*(19)+in_buf[43]*(0)+in_buf[44]*(13)+in_buf[45]*(-8)+in_buf[46]*(-19)+in_buf[47]*(-22)+in_buf[48]*(-20)+in_buf[49]*(-25)+in_buf[50]*(-17)+in_buf[51]*(-9)+in_buf[52]*(3)+in_buf[53]*(2)+in_buf[54]*(3)+in_buf[55]*(-3)+in_buf[56]*(1)+in_buf[57]*(-3)+in_buf[58]*(-11)+in_buf[59]*(-30)+in_buf[60]*(-38)+in_buf[61]*(-8)+in_buf[62]*(-7)+in_buf[63]*(-20)+in_buf[64]*(-21)+in_buf[65]*(-24)+in_buf[66]*(-27)+in_buf[67]*(-25)+in_buf[68]*(-39)+in_buf[69]*(-15)+in_buf[70]*(3)+in_buf[71]*(16)+in_buf[72]*(15)+in_buf[73]*(14)+in_buf[74]*(0)+in_buf[75]*(-9)+in_buf[76]*(2)+in_buf[77]*(9)+in_buf[78]*(-16)+in_buf[79]*(-15)+in_buf[80]*(12)+in_buf[81]*(-1)+in_buf[82]*(3)+in_buf[83]*(-2)+in_buf[84]*(0)+in_buf[85]*(-1)+in_buf[86]*(0)+in_buf[87]*(-35)+in_buf[88]*(-39)+in_buf[89]*(-25)+in_buf[90]*(-31)+in_buf[91]*(-21)+in_buf[92]*(-35)+in_buf[93]*(-23)+in_buf[94]*(-4)+in_buf[95]*(19)+in_buf[96]*(-18)+in_buf[97]*(-9)+in_buf[98]*(18)+in_buf[99]*(22)+in_buf[100]*(29)+in_buf[101]*(22)+in_buf[102]*(18)+in_buf[103]*(10)+in_buf[104]*(11)+in_buf[105]*(2)+in_buf[106]*(-2)+in_buf[107]*(-24)+in_buf[108]*(-31)+in_buf[109]*(11)+in_buf[110]*(-23)+in_buf[111]*(-3)+in_buf[112]*(0)+in_buf[113]*(5)+in_buf[114]*(10)+in_buf[115]*(-9)+in_buf[116]*(-29)+in_buf[117]*(-24)+in_buf[118]*(-22)+in_buf[119]*(-10)+in_buf[120]*(-15)+in_buf[121]*(5)+in_buf[122]*(10)+in_buf[123]*(0)+in_buf[124]*(5)+in_buf[125]*(3)+in_buf[126]*(-3)+in_buf[127]*(7)+in_buf[128]*(14)+in_buf[129]*(23)+in_buf[130]*(29)+in_buf[131]*(19)+in_buf[132]*(17)+in_buf[133]*(-6)+in_buf[134]*(17)+in_buf[135]*(-13)+in_buf[136]*(-18)+in_buf[137]*(-9)+in_buf[138]*(-35)+in_buf[139]*(-22)+in_buf[140]*(2)+in_buf[141]*(0)+in_buf[142]*(-4)+in_buf[143]*(-2)+in_buf[144]*(-26)+in_buf[145]*(-9)+in_buf[146]*(-15)+in_buf[147]*(-2)+in_buf[148]*(4)+in_buf[149]*(-5)+in_buf[150]*(-18)+in_buf[151]*(-35)+in_buf[152]*(-13)+in_buf[153]*(-17)+in_buf[154]*(-13)+in_buf[155]*(0)+in_buf[156]*(8)+in_buf[157]*(12)+in_buf[158]*(32)+in_buf[159]*(36)+in_buf[160]*(20)+in_buf[161]*(-5)+in_buf[162]*(17)+in_buf[163]*(27)+in_buf[164]*(5)+in_buf[165]*(27)+in_buf[166]*(-47)+in_buf[167]*(-24)+in_buf[168]*(0)+in_buf[169]*(16)+in_buf[170]*(-8)+in_buf[171]*(3)+in_buf[172]*(7)+in_buf[173]*(-19)+in_buf[174]*(-3)+in_buf[175]*(-1)+in_buf[176]*(-5)+in_buf[177]*(0)+in_buf[178]*(-16)+in_buf[179]*(-21)+in_buf[180]*(-4)+in_buf[181]*(-10)+in_buf[182]*(-18)+in_buf[183]*(-25)+in_buf[184]*(-3)+in_buf[185]*(19)+in_buf[186]*(29)+in_buf[187]*(37)+in_buf[188]*(27)+in_buf[189]*(-2)+in_buf[190]*(-9)+in_buf[191]*(3)+in_buf[192]*(-20)+in_buf[193]*(-24)+in_buf[194]*(-5)+in_buf[195]*(-20)+in_buf[196]*(0)+in_buf[197]*(32)+in_buf[198]*(4)+in_buf[199]*(30)+in_buf[200]*(15)+in_buf[201]*(-21)+in_buf[202]*(-1)+in_buf[203]*(5)+in_buf[204]*(-13)+in_buf[205]*(-17)+in_buf[206]*(-4)+in_buf[207]*(-3)+in_buf[208]*(3)+in_buf[209]*(-2)+in_buf[210]*(-27)+in_buf[211]*(-37)+in_buf[212]*(-20)+in_buf[213]*(14)+in_buf[214]*(32)+in_buf[215]*(45)+in_buf[216]*(41)+in_buf[217]*(18)+in_buf[218]*(5)+in_buf[219]*(4)+in_buf[220]*(-3)+in_buf[221]*(-46)+in_buf[222]*(-34)+in_buf[223]*(-24)+in_buf[224]*(-20)+in_buf[225]*(21)+in_buf[226]*(34)+in_buf[227]*(11)+in_buf[228]*(-18)+in_buf[229]*(-22)+in_buf[230]*(-3)+in_buf[231]*(11)+in_buf[232]*(-5)+in_buf[233]*(-13)+in_buf[234]*(3)+in_buf[235]*(0)+in_buf[236]*(-13)+in_buf[237]*(-8)+in_buf[238]*(-36)+in_buf[239]*(-40)+in_buf[240]*(-33)+in_buf[241]*(12)+in_buf[242]*(48)+in_buf[243]*(51)+in_buf[244]*(30)+in_buf[245]*(24)+in_buf[246]*(18)+in_buf[247]*(6)+in_buf[248]*(-21)+in_buf[249]*(-18)+in_buf[250]*(-11)+in_buf[251]*(-9)+in_buf[252]*(6)+in_buf[253]*(14)+in_buf[254]*(17)+in_buf[255]*(16)+in_buf[256]*(-10)+in_buf[257]*(-6)+in_buf[258]*(3)+in_buf[259]*(1)+in_buf[260]*(3)+in_buf[261]*(6)+in_buf[262]*(10)+in_buf[263]*(-12)+in_buf[264]*(-5)+in_buf[265]*(-15)+in_buf[266]*(-50)+in_buf[267]*(-58)+in_buf[268]*(-20)+in_buf[269]*(23)+in_buf[270]*(55)+in_buf[271]*(50)+in_buf[272]*(33)+in_buf[273]*(28)+in_buf[274]*(20)+in_buf[275]*(6)+in_buf[276]*(-39)+in_buf[277]*(-15)+in_buf[278]*(-27)+in_buf[279]*(-4)+in_buf[280]*(17)+in_buf[281]*(8)+in_buf[282]*(7)+in_buf[283]*(3)+in_buf[284]*(-16)+in_buf[285]*(-4)+in_buf[286]*(0)+in_buf[287]*(0)+in_buf[288]*(10)+in_buf[289]*(11)+in_buf[290]*(-6)+in_buf[291]*(-2)+in_buf[292]*(-12)+in_buf[293]*(-20)+in_buf[294]*(-49)+in_buf[295]*(-68)+in_buf[296]*(-24)+in_buf[297]*(44)+in_buf[298]*(45)+in_buf[299]*(52)+in_buf[300]*(30)+in_buf[301]*(25)+in_buf[302]*(21)+in_buf[303]*(-11)+in_buf[304]*(-38)+in_buf[305]*(-14)+in_buf[306]*(-48)+in_buf[307]*(-3)+in_buf[308]*(17)+in_buf[309]*(-29)+in_buf[310]*(-39)+in_buf[311]*(-14)+in_buf[312]*(-20)+in_buf[313]*(4)+in_buf[314]*(2)+in_buf[315]*(-3)+in_buf[316]*(6)+in_buf[317]*(-7)+in_buf[318]*(-9)+in_buf[319]*(-17)+in_buf[320]*(-18)+in_buf[321]*(-12)+in_buf[322]*(-46)+in_buf[323]*(-38)+in_buf[324]*(-1)+in_buf[325]*(28)+in_buf[326]*(32)+in_buf[327]*(36)+in_buf[328]*(32)+in_buf[329]*(14)+in_buf[330]*(3)+in_buf[331]*(-19)+in_buf[332]*(-20)+in_buf[333]*(5)+in_buf[334]*(-37)+in_buf[335]*(-5)+in_buf[336]*(13)+in_buf[337]*(-2)+in_buf[338]*(-25)+in_buf[339]*(-15)+in_buf[340]*(0)+in_buf[341]*(0)+in_buf[342]*(2)+in_buf[343]*(-17)+in_buf[344]*(-5)+in_buf[345]*(-18)+in_buf[346]*(-11)+in_buf[347]*(-21)+in_buf[348]*(-3)+in_buf[349]*(-16)+in_buf[350]*(-25)+in_buf[351]*(-19)+in_buf[352]*(-3)+in_buf[353]*(25)+in_buf[354]*(22)+in_buf[355]*(21)+in_buf[356]*(-1)+in_buf[357]*(-1)+in_buf[358]*(-8)+in_buf[359]*(-18)+in_buf[360]*(-6)+in_buf[361]*(-2)+in_buf[362]*(-14)+in_buf[363]*(-5)+in_buf[364]*(-4)+in_buf[365]*(-5)+in_buf[366]*(13)+in_buf[367]*(-23)+in_buf[368]*(1)+in_buf[369]*(6)+in_buf[370]*(3)+in_buf[371]*(-24)+in_buf[372]*(1)+in_buf[373]*(-8)+in_buf[374]*(-8)+in_buf[375]*(-5)+in_buf[376]*(-14)+in_buf[377]*(-18)+in_buf[378]*(-14)+in_buf[379]*(-13)+in_buf[380]*(-3)+in_buf[381]*(23)+in_buf[382]*(19)+in_buf[383]*(3)+in_buf[384]*(0)+in_buf[385]*(-1)+in_buf[386]*(-3)+in_buf[387]*(-17)+in_buf[388]*(1)+in_buf[389]*(11)+in_buf[390]*(4)+in_buf[391]*(-5)+in_buf[392]*(-1)+in_buf[393]*(5)+in_buf[394]*(0)+in_buf[395]*(-26)+in_buf[396]*(8)+in_buf[397]*(0)+in_buf[398]*(15)+in_buf[399]*(18)+in_buf[400]*(5)+in_buf[401]*(2)+in_buf[402]*(-2)+in_buf[403]*(-3)+in_buf[404]*(1)+in_buf[405]*(-9)+in_buf[406]*(-1)+in_buf[407]*(3)+in_buf[408]*(19)+in_buf[409]*(28)+in_buf[410]*(8)+in_buf[411]*(14)+in_buf[412]*(2)+in_buf[413]*(-19)+in_buf[414]*(-9)+in_buf[415]*(-34)+in_buf[416]*(-12)+in_buf[417]*(15)+in_buf[418]*(15)+in_buf[419]*(4)+in_buf[420]*(5)+in_buf[421]*(5)+in_buf[422]*(12)+in_buf[423]*(10)+in_buf[424]*(22)+in_buf[425]*(15)+in_buf[426]*(2)+in_buf[427]*(8)+in_buf[428]*(12)+in_buf[429]*(2)+in_buf[430]*(0)+in_buf[431]*(-4)+in_buf[432]*(-9)+in_buf[433]*(-2)+in_buf[434]*(-3)+in_buf[435]*(11)+in_buf[436]*(11)+in_buf[437]*(15)+in_buf[438]*(14)+in_buf[439]*(15)+in_buf[440]*(0)+in_buf[441]*(-13)+in_buf[442]*(6)+in_buf[443]*(-12)+in_buf[444]*(-18)+in_buf[445]*(16)+in_buf[446]*(39)+in_buf[447]*(4)+in_buf[448]*(6)+in_buf[449]*(15)+in_buf[450]*(14)+in_buf[451]*(-13)+in_buf[452]*(14)+in_buf[453]*(24)+in_buf[454]*(3)+in_buf[455]*(0)+in_buf[456]*(-7)+in_buf[457]*(-2)+in_buf[458]*(-2)+in_buf[459]*(-17)+in_buf[460]*(-4)+in_buf[461]*(0)+in_buf[462]*(2)+in_buf[463]*(6)+in_buf[464]*(6)+in_buf[465]*(15)+in_buf[466]*(2)+in_buf[467]*(9)+in_buf[468]*(2)+in_buf[469]*(2)+in_buf[470]*(0)+in_buf[471]*(11)+in_buf[472]*(12)+in_buf[473]*(16)+in_buf[474]*(38)+in_buf[475]*(9)+in_buf[476]*(1)+in_buf[477]*(6)+in_buf[478]*(31)+in_buf[479]*(1)+in_buf[480]*(15)+in_buf[481]*(14)+in_buf[482]*(5)+in_buf[483]*(4)+in_buf[484]*(-6)+in_buf[485]*(-13)+in_buf[486]*(-11)+in_buf[487]*(-8)+in_buf[488]*(-1)+in_buf[489]*(3)+in_buf[490]*(-8)+in_buf[491]*(1)+in_buf[492]*(4)+in_buf[493]*(7)+in_buf[494]*(0)+in_buf[495]*(3)+in_buf[496]*(-7)+in_buf[497]*(0)+in_buf[498]*(-9)+in_buf[499]*(7)+in_buf[500]*(15)+in_buf[501]*(37)+in_buf[502]*(41)+in_buf[503]*(2)+in_buf[504]*(10)+in_buf[505]*(13)+in_buf[506]*(30)+in_buf[507]*(4)+in_buf[508]*(9)+in_buf[509]*(8)+in_buf[510]*(1)+in_buf[511]*(5)+in_buf[512]*(-3)+in_buf[513]*(-7)+in_buf[514]*(-26)+in_buf[515]*(-12)+in_buf[516]*(-11)+in_buf[517]*(5)+in_buf[518]*(4)+in_buf[519]*(6)+in_buf[520]*(16)+in_buf[521]*(12)+in_buf[522]*(15)+in_buf[523]*(0)+in_buf[524]*(-10)+in_buf[525]*(-10)+in_buf[526]*(-1)+in_buf[527]*(7)+in_buf[528]*(7)+in_buf[529]*(8)+in_buf[530]*(14)+in_buf[531]*(0)+in_buf[532]*(2)+in_buf[533]*(-11)+in_buf[534]*(-6)+in_buf[535]*(3)+in_buf[536]*(9)+in_buf[537]*(14)+in_buf[538]*(8)+in_buf[539]*(19)+in_buf[540]*(6)+in_buf[541]*(7)+in_buf[542]*(-6)+in_buf[543]*(-9)+in_buf[544]*(-13)+in_buf[545]*(8)+in_buf[546]*(-2)+in_buf[547]*(8)+in_buf[548]*(19)+in_buf[549]*(20)+in_buf[550]*(-3)+in_buf[551]*(3)+in_buf[552]*(-15)+in_buf[553]*(2)+in_buf[554]*(2)+in_buf[555]*(0)+in_buf[556]*(-6)+in_buf[557]*(-2)+in_buf[558]*(20)+in_buf[559]*(5)+in_buf[560]*(-1)+in_buf[561]*(-10)+in_buf[562]*(5)+in_buf[563]*(14)+in_buf[564]*(1)+in_buf[565]*(11)+in_buf[566]*(12)+in_buf[567]*(14)+in_buf[568]*(0)+in_buf[569]*(-1)+in_buf[570]*(5)+in_buf[571]*(4)+in_buf[572]*(1)+in_buf[573]*(-6)+in_buf[574]*(-8)+in_buf[575]*(-1)+in_buf[576]*(12)+in_buf[577]*(11)+in_buf[578]*(5)+in_buf[579]*(8)+in_buf[580]*(9)+in_buf[581]*(12)+in_buf[582]*(-4)+in_buf[583]*(2)+in_buf[584]*(9)+in_buf[585]*(-14)+in_buf[586]*(20)+in_buf[587]*(7)+in_buf[588]*(-1)+in_buf[589]*(2)+in_buf[590]*(41)+in_buf[591]*(24)+in_buf[592]*(0)+in_buf[593]*(5)+in_buf[594]*(12)+in_buf[595]*(5)+in_buf[596]*(8)+in_buf[597]*(5)+in_buf[598]*(23)+in_buf[599]*(7)+in_buf[600]*(0)+in_buf[601]*(-11)+in_buf[602]*(-22)+in_buf[603]*(-11)+in_buf[604]*(15)+in_buf[605]*(17)+in_buf[606]*(17)+in_buf[607]*(10)+in_buf[608]*(13)+in_buf[609]*(10)+in_buf[610]*(13)+in_buf[611]*(0)+in_buf[612]*(17)+in_buf[613]*(-8)+in_buf[614]*(-24)+in_buf[615]*(3)+in_buf[616]*(-2)+in_buf[617]*(-1)+in_buf[618]*(41)+in_buf[619]*(-16)+in_buf[620]*(-10)+in_buf[621]*(-2)+in_buf[622]*(8)+in_buf[623]*(16)+in_buf[624]*(18)+in_buf[625]*(5)+in_buf[626]*(8)+in_buf[627]*(10)+in_buf[628]*(0)+in_buf[629]*(-15)+in_buf[630]*(-17)+in_buf[631]*(-2)+in_buf[632]*(-2)+in_buf[633]*(8)+in_buf[634]*(4)+in_buf[635]*(10)+in_buf[636]*(-1)+in_buf[637]*(13)+in_buf[638]*(25)+in_buf[639]*(2)+in_buf[640]*(20)+in_buf[641]*(-1)+in_buf[642]*(-12)+in_buf[643]*(4)+in_buf[644]*(0)+in_buf[645]*(2)+in_buf[646]*(8)+in_buf[647]*(-34)+in_buf[648]*(-36)+in_buf[649]*(-13)+in_buf[650]*(9)+in_buf[651]*(24)+in_buf[652]*(5)+in_buf[653]*(1)+in_buf[654]*(16)+in_buf[655]*(15)+in_buf[656]*(-8)+in_buf[657]*(-26)+in_buf[658]*(-18)+in_buf[659]*(2)+in_buf[660]*(0)+in_buf[661]*(-17)+in_buf[662]*(-3)+in_buf[663]*(6)+in_buf[664]*(2)+in_buf[665]*(21)+in_buf[666]*(18)+in_buf[667]*(16)+in_buf[668]*(16)+in_buf[669]*(0)+in_buf[670]*(-16)+in_buf[671]*(0)+in_buf[672]*(4)+in_buf[673]*(4)+in_buf[674]*(17)+in_buf[675]*(-9)+in_buf[676]*(18)+in_buf[677]*(-18)+in_buf[678]*(11)+in_buf[679]*(18)+in_buf[680]*(13)+in_buf[681]*(5)+in_buf[682]*(14)+in_buf[683]*(15)+in_buf[684]*(3)+in_buf[685]*(-25)+in_buf[686]*(-18)+in_buf[687]*(-19)+in_buf[688]*(-10)+in_buf[689]*(-7)+in_buf[690]*(-14)+in_buf[691]*(-22)+in_buf[692]*(-12)+in_buf[693]*(19)+in_buf[694]*(19)+in_buf[695]*(21)+in_buf[696]*(12)+in_buf[697]*(19)+in_buf[698]*(17)+in_buf[699]*(3)+in_buf[700]*(2)+in_buf[701]*(0)+in_buf[702]*(-20)+in_buf[703]*(12)+in_buf[704]*(5)+in_buf[705]*(-6)+in_buf[706]*(9)+in_buf[707]*(8)+in_buf[708]*(28)+in_buf[709]*(20)+in_buf[710]*(9)+in_buf[711]*(4)+in_buf[712]*(5)+in_buf[713]*(-13)+in_buf[714]*(14)+in_buf[715]*(3)+in_buf[716]*(16)+in_buf[717]*(0)+in_buf[718]*(8)+in_buf[719]*(-27)+in_buf[720]*(-19)+in_buf[721]*(-15)+in_buf[722]*(-31)+in_buf[723]*(-17)+in_buf[724]*(-27)+in_buf[725]*(1)+in_buf[726]*(8)+in_buf[727]*(0)+in_buf[728]*(-3)+in_buf[729]*(2)+in_buf[730]*(3)+in_buf[731]*(3)+in_buf[732]*(-8)+in_buf[733]*(-26)+in_buf[734]*(14)+in_buf[735]*(23)+in_buf[736]*(-6)+in_buf[737]*(4)+in_buf[738]*(-3)+in_buf[739]*(-22)+in_buf[740]*(-15)+in_buf[741]*(2)+in_buf[742]*(18)+in_buf[743]*(20)+in_buf[744]*(-1)+in_buf[745]*(-4)+in_buf[746]*(-11)+in_buf[747]*(-36)+in_buf[748]*(-6)+in_buf[749]*(9)+in_buf[750]*(-9)+in_buf[751]*(15)+in_buf[752]*(19)+in_buf[753]*(6)+in_buf[754]*(0)+in_buf[755]*(3)+in_buf[756]*(-3)+in_buf[757]*(1)+in_buf[758]*(-3)+in_buf[759]*(-1)+in_buf[760]*(25)+in_buf[761]*(26)+in_buf[762]*(24)+in_buf[763]*(0)+in_buf[764]*(-7)+in_buf[765]*(0)+in_buf[766]*(-22)+in_buf[767]*(-3)+in_buf[768]*(-4)+in_buf[769]*(44)+in_buf[770]*(39)+in_buf[771]*(34)+in_buf[772]*(8)+in_buf[773]*(32)+in_buf[774]*(23)+in_buf[775]*(-9)+in_buf[776]*(13)+in_buf[777]*(35)+in_buf[778]*(-2)+in_buf[779]*(18)+in_buf[780]*(-3)+in_buf[781]*(-2)+in_buf[782]*(2)+in_buf[783]*(2);
assign in_buf_weight032=in_buf[0]*(1)+in_buf[1]*(4)+in_buf[2]*(0)+in_buf[3]*(-2)+in_buf[4]*(4)+in_buf[5]*(0)+in_buf[6]*(-2)+in_buf[7]*(1)+in_buf[8]*(1)+in_buf[9]*(-2)+in_buf[10]*(-2)+in_buf[11]*(4)+in_buf[12]*(4)+in_buf[13]*(1)+in_buf[14]*(-4)+in_buf[15]*(-2)+in_buf[16]*(-1)+in_buf[17]*(-1)+in_buf[18]*(2)+in_buf[19]*(1)+in_buf[20]*(-2)+in_buf[21]*(3)+in_buf[22]*(1)+in_buf[23]*(2)+in_buf[24]*(2)+in_buf[25]*(-3)+in_buf[26]*(-3)+in_buf[27]*(-3)+in_buf[28]*(-3)+in_buf[29]*(-3)+in_buf[30]*(3)+in_buf[31]*(-1)+in_buf[32]*(6)+in_buf[33]*(-8)+in_buf[34]*(-4)+in_buf[35]*(-8)+in_buf[36]*(-3)+in_buf[37]*(5)+in_buf[38]*(8)+in_buf[39]*(6)+in_buf[40]*(3)+in_buf[41]*(24)+in_buf[42]*(20)+in_buf[43]*(-29)+in_buf[44]*(-29)+in_buf[45]*(-22)+in_buf[46]*(3)+in_buf[47]*(0)+in_buf[48]*(8)+in_buf[49]*(18)+in_buf[50]*(11)+in_buf[51]*(-3)+in_buf[52]*(3)+in_buf[53]*(-1)+in_buf[54]*(0)+in_buf[55]*(2)+in_buf[56]*(0)+in_buf[57]*(-3)+in_buf[58]*(2)+in_buf[59]*(-7)+in_buf[60]*(-4)+in_buf[61]*(-1)+in_buf[62]*(0)+in_buf[63]*(-12)+in_buf[64]*(2)+in_buf[65]*(-1)+in_buf[66]*(-6)+in_buf[67]*(16)+in_buf[68]*(-3)+in_buf[69]*(-4)+in_buf[70]*(31)+in_buf[71]*(16)+in_buf[72]*(-37)+in_buf[73]*(-12)+in_buf[74]*(3)+in_buf[75]*(3)+in_buf[76]*(-4)+in_buf[77]*(-13)+in_buf[78]*(0)+in_buf[79]*(-12)+in_buf[80]*(-10)+in_buf[81]*(-8)+in_buf[82]*(1)+in_buf[83]*(4)+in_buf[84]*(-3)+in_buf[85]*(-1)+in_buf[86]*(-3)+in_buf[87]*(-9)+in_buf[88]*(-4)+in_buf[89]*(13)+in_buf[90]*(7)+in_buf[91]*(6)+in_buf[92]*(4)+in_buf[93]*(-34)+in_buf[94]*(-18)+in_buf[95]*(2)+in_buf[96]*(2)+in_buf[97]*(-8)+in_buf[98]*(-12)+in_buf[99]*(-12)+in_buf[100]*(-15)+in_buf[101]*(-19)+in_buf[102]*(-13)+in_buf[103]*(9)+in_buf[104]*(36)+in_buf[105]*(54)+in_buf[106]*(23)+in_buf[107]*(-1)+in_buf[108]*(-11)+in_buf[109]*(-12)+in_buf[110]*(1)+in_buf[111]*(4)+in_buf[112]*(0)+in_buf[113]*(-6)+in_buf[114]*(2)+in_buf[115]*(14)+in_buf[116]*(3)+in_buf[117]*(-34)+in_buf[118]*(-30)+in_buf[119]*(11)+in_buf[120]*(-15)+in_buf[121]*(-4)+in_buf[122]*(5)+in_buf[123]*(22)+in_buf[124]*(24)+in_buf[125]*(6)+in_buf[126]*(14)+in_buf[127]*(3)+in_buf[128]*(17)+in_buf[129]*(12)+in_buf[130]*(-11)+in_buf[131]*(0)+in_buf[132]*(4)+in_buf[133]*(0)+in_buf[134]*(-3)+in_buf[135]*(33)+in_buf[136]*(52)+in_buf[137]*(48)+in_buf[138]*(71)+in_buf[139]*(29)+in_buf[140]*(0)+in_buf[141]*(-1)+in_buf[142]*(-5)+in_buf[143]*(-21)+in_buf[144]*(-27)+in_buf[145]*(-29)+in_buf[146]*(5)+in_buf[147]*(15)+in_buf[148]*(24)+in_buf[149]*(40)+in_buf[150]*(18)+in_buf[151]*(24)+in_buf[152]*(8)+in_buf[153]*(-7)+in_buf[154]*(1)+in_buf[155]*(-11)+in_buf[156]*(-2)+in_buf[157]*(5)+in_buf[158]*(-17)+in_buf[159]*(-21)+in_buf[160]*(-4)+in_buf[161]*(0)+in_buf[162]*(0)+in_buf[163]*(0)+in_buf[164]*(23)+in_buf[165]*(52)+in_buf[166]*(48)+in_buf[167]*(28)+in_buf[168]*(1)+in_buf[169]*(-1)+in_buf[170]*(20)+in_buf[171]*(-55)+in_buf[172]*(-10)+in_buf[173]*(22)+in_buf[174]*(7)+in_buf[175]*(26)+in_buf[176]*(31)+in_buf[177]*(23)+in_buf[178]*(3)+in_buf[179]*(1)+in_buf[180]*(-3)+in_buf[181]*(-6)+in_buf[182]*(-8)+in_buf[183]*(-7)+in_buf[184]*(-16)+in_buf[185]*(0)+in_buf[186]*(-5)+in_buf[187]*(-2)+in_buf[188]*(-12)+in_buf[189]*(-9)+in_buf[190]*(13)+in_buf[191]*(13)+in_buf[192]*(25)+in_buf[193]*(70)+in_buf[194]*(24)+in_buf[195]*(-19)+in_buf[196]*(-1)+in_buf[197]*(-24)+in_buf[198]*(11)+in_buf[199]*(-56)+in_buf[200]*(-21)+in_buf[201]*(23)+in_buf[202]*(14)+in_buf[203]*(17)+in_buf[204]*(30)+in_buf[205]*(17)+in_buf[206]*(8)+in_buf[207]*(-7)+in_buf[208]*(-15)+in_buf[209]*(-22)+in_buf[210]*(-26)+in_buf[211]*(-9)+in_buf[212]*(-1)+in_buf[213]*(-1)+in_buf[214]*(11)+in_buf[215]*(15)+in_buf[216]*(4)+in_buf[217]*(1)+in_buf[218]*(8)+in_buf[219]*(14)+in_buf[220]*(34)+in_buf[221]*(45)+in_buf[222]*(27)+in_buf[223]*(-12)+in_buf[224]*(-2)+in_buf[225]*(-33)+in_buf[226]*(10)+in_buf[227]*(4)+in_buf[228]*(3)+in_buf[229]*(26)+in_buf[230]*(28)+in_buf[231]*(32)+in_buf[232]*(26)+in_buf[233]*(24)+in_buf[234]*(-3)+in_buf[235]*(-2)+in_buf[236]*(-11)+in_buf[237]*(-28)+in_buf[238]*(-33)+in_buf[239]*(-10)+in_buf[240]*(9)+in_buf[241]*(8)+in_buf[242]*(7)+in_buf[243]*(5)+in_buf[244]*(11)+in_buf[245]*(10)+in_buf[246]*(7)+in_buf[247]*(25)+in_buf[248]*(54)+in_buf[249]*(56)+in_buf[250]*(33)+in_buf[251]*(37)+in_buf[252]*(-1)+in_buf[253]*(-14)+in_buf[254]*(-3)+in_buf[255]*(-7)+in_buf[256]*(-3)+in_buf[257]*(1)+in_buf[258]*(29)+in_buf[259]*(15)+in_buf[260]*(17)+in_buf[261]*(18)+in_buf[262]*(13)+in_buf[263]*(17)+in_buf[264]*(-19)+in_buf[265]*(-42)+in_buf[266]*(-33)+in_buf[267]*(-5)+in_buf[268]*(16)+in_buf[269]*(-1)+in_buf[270]*(-4)+in_buf[271]*(-4)+in_buf[272]*(13)+in_buf[273]*(20)+in_buf[274]*(19)+in_buf[275]*(33)+in_buf[276]*(34)+in_buf[277]*(40)+in_buf[278]*(10)+in_buf[279]*(-20)+in_buf[280]*(-2)+in_buf[281]*(-5)+in_buf[282]*(-35)+in_buf[283]*(-14)+in_buf[284]*(25)+in_buf[285]*(11)+in_buf[286]*(10)+in_buf[287]*(16)+in_buf[288]*(16)+in_buf[289]*(34)+in_buf[290]*(36)+in_buf[291]*(27)+in_buf[292]*(4)+in_buf[293]*(-42)+in_buf[294]*(-40)+in_buf[295]*(-9)+in_buf[296]*(-19)+in_buf[297]*(-24)+in_buf[298]*(-9)+in_buf[299]*(-5)+in_buf[300]*(1)+in_buf[301]*(0)+in_buf[302]*(20)+in_buf[303]*(23)+in_buf[304]*(19)+in_buf[305]*(0)+in_buf[306]*(11)+in_buf[307]*(-10)+in_buf[308]*(6)+in_buf[309]*(-40)+in_buf[310]*(-26)+in_buf[311]*(-6)+in_buf[312]*(16)+in_buf[313]*(17)+in_buf[314]*(11)+in_buf[315]*(12)+in_buf[316]*(34)+in_buf[317]*(43)+in_buf[318]*(37)+in_buf[319]*(43)+in_buf[320]*(27)+in_buf[321]*(-16)+in_buf[322]*(-16)+in_buf[323]*(-11)+in_buf[324]*(-25)+in_buf[325]*(-25)+in_buf[326]*(-24)+in_buf[327]*(-13)+in_buf[328]*(-7)+in_buf[329]*(-1)+in_buf[330]*(2)+in_buf[331]*(-5)+in_buf[332]*(1)+in_buf[333]*(0)+in_buf[334]*(45)+in_buf[335]*(-16)+in_buf[336]*(9)+in_buf[337]*(-2)+in_buf[338]*(-13)+in_buf[339]*(4)+in_buf[340]*(-4)+in_buf[341]*(0)+in_buf[342]*(14)+in_buf[343]*(28)+in_buf[344]*(30)+in_buf[345]*(36)+in_buf[346]*(40)+in_buf[347]*(35)+in_buf[348]*(33)+in_buf[349]*(9)+in_buf[350]*(-22)+in_buf[351]*(-11)+in_buf[352]*(-9)+in_buf[353]*(-13)+in_buf[354]*(-7)+in_buf[355]*(1)+in_buf[356]*(2)+in_buf[357]*(8)+in_buf[358]*(2)+in_buf[359]*(7)+in_buf[360]*(12)+in_buf[361]*(-1)+in_buf[362]*(9)+in_buf[363]*(-30)+in_buf[364]*(1)+in_buf[365]*(4)+in_buf[366]*(-16)+in_buf[367]*(0)+in_buf[368]*(-14)+in_buf[369]*(21)+in_buf[370]*(8)+in_buf[371]*(19)+in_buf[372]*(22)+in_buf[373]*(29)+in_buf[374]*(28)+in_buf[375]*(37)+in_buf[376]*(32)+in_buf[377]*(11)+in_buf[378]*(-6)+in_buf[379]*(16)+in_buf[380]*(8)+in_buf[381]*(-7)+in_buf[382]*(4)+in_buf[383]*(7)+in_buf[384]*(9)+in_buf[385]*(-4)+in_buf[386]*(13)+in_buf[387]*(10)+in_buf[388]*(4)+in_buf[389]*(-10)+in_buf[390]*(-11)+in_buf[391]*(-12)+in_buf[392]*(21)+in_buf[393]*(-6)+in_buf[394]*(-18)+in_buf[395]*(3)+in_buf[396]*(-6)+in_buf[397]*(34)+in_buf[398]*(17)+in_buf[399]*(9)+in_buf[400]*(21)+in_buf[401]*(15)+in_buf[402]*(22)+in_buf[403]*(38)+in_buf[404]*(21)+in_buf[405]*(6)+in_buf[406]*(12)+in_buf[407]*(7)+in_buf[408]*(6)+in_buf[409]*(19)+in_buf[410]*(0)+in_buf[411]*(6)+in_buf[412]*(-10)+in_buf[413]*(-10)+in_buf[414]*(4)+in_buf[415]*(7)+in_buf[416]*(6)+in_buf[417]*(-24)+in_buf[418]*(-35)+in_buf[419]*(-18)+in_buf[420]*(16)+in_buf[421]*(5)+in_buf[422]*(23)+in_buf[423]*(2)+in_buf[424]*(7)+in_buf[425]*(2)+in_buf[426]*(11)+in_buf[427]*(1)+in_buf[428]*(0)+in_buf[429]*(19)+in_buf[430]*(15)+in_buf[431]*(25)+in_buf[432]*(24)+in_buf[433]*(15)+in_buf[434]*(16)+in_buf[435]*(10)+in_buf[436]*(3)+in_buf[437]*(17)+in_buf[438]*(-5)+in_buf[439]*(-7)+in_buf[440]*(-14)+in_buf[441]*(-25)+in_buf[442]*(-5)+in_buf[443]*(18)+in_buf[444]*(0)+in_buf[445]*(3)+in_buf[446]*(10)+in_buf[447]*(-14)+in_buf[448]*(-8)+in_buf[449]*(0)+in_buf[450]*(8)+in_buf[451]*(-12)+in_buf[452]*(-42)+in_buf[453]*(-17)+in_buf[454]*(-14)+in_buf[455]*(-23)+in_buf[456]*(-12)+in_buf[457]*(-2)+in_buf[458]*(1)+in_buf[459]*(4)+in_buf[460]*(23)+in_buf[461]*(30)+in_buf[462]*(12)+in_buf[463]*(13)+in_buf[464]*(10)+in_buf[465]*(3)+in_buf[466]*(-2)+in_buf[467]*(-5)+in_buf[468]*(-5)+in_buf[469]*(-13)+in_buf[470]*(0)+in_buf[471]*(9)+in_buf[472]*(-15)+in_buf[473]*(6)+in_buf[474]*(-18)+in_buf[475]*(-20)+in_buf[476]*(2)+in_buf[477]*(1)+in_buf[478]*(4)+in_buf[479]*(-1)+in_buf[480]*(-34)+in_buf[481]*(-21)+in_buf[482]*(-24)+in_buf[483]*(-38)+in_buf[484]*(-26)+in_buf[485]*(-7)+in_buf[486]*(0)+in_buf[487]*(12)+in_buf[488]*(24)+in_buf[489]*(20)+in_buf[490]*(-2)+in_buf[491]*(-3)+in_buf[492]*(9)+in_buf[493]*(-5)+in_buf[494]*(-1)+in_buf[495]*(-3)+in_buf[496]*(16)+in_buf[497]*(10)+in_buf[498]*(-2)+in_buf[499]*(6)+in_buf[500]*(0)+in_buf[501]*(-30)+in_buf[502]*(-15)+in_buf[503]*(-18)+in_buf[504]*(-29)+in_buf[505]*(-3)+in_buf[506]*(-7)+in_buf[507]*(-1)+in_buf[508]*(-31)+in_buf[509]*(4)+in_buf[510]*(-14)+in_buf[511]*(-54)+in_buf[512]*(-36)+in_buf[513]*(-17)+in_buf[514]*(-3)+in_buf[515]*(2)+in_buf[516]*(16)+in_buf[517]*(11)+in_buf[518]*(-12)+in_buf[519]*(-16)+in_buf[520]*(-1)+in_buf[521]*(-11)+in_buf[522]*(-15)+in_buf[523]*(-1)+in_buf[524]*(9)+in_buf[525]*(-7)+in_buf[526]*(-18)+in_buf[527]*(-8)+in_buf[528]*(-10)+in_buf[529]*(-65)+in_buf[530]*(-25)+in_buf[531]*(-3)+in_buf[532]*(1)+in_buf[533]*(-32)+in_buf[534]*(-43)+in_buf[535]*(-7)+in_buf[536]*(-36)+in_buf[537]*(12)+in_buf[538]*(-6)+in_buf[539]*(-36)+in_buf[540]*(-10)+in_buf[541]*(-16)+in_buf[542]*(-13)+in_buf[543]*(-11)+in_buf[544]*(6)+in_buf[545]*(-4)+in_buf[546]*(-7)+in_buf[547]*(-9)+in_buf[548]*(-11)+in_buf[549]*(-11)+in_buf[550]*(-11)+in_buf[551]*(-7)+in_buf[552]*(0)+in_buf[553]*(-9)+in_buf[554]*(1)+in_buf[555]*(13)+in_buf[556]*(1)+in_buf[557]*(-42)+in_buf[558]*(-30)+in_buf[559]*(-5)+in_buf[560]*(3)+in_buf[561]*(-2)+in_buf[562]*(-17)+in_buf[563]*(-39)+in_buf[564]*(-45)+in_buf[565]*(-11)+in_buf[566]*(-23)+in_buf[567]*(-20)+in_buf[568]*(0)+in_buf[569]*(0)+in_buf[570]*(-4)+in_buf[571]*(-13)+in_buf[572]*(-4)+in_buf[573]*(-9)+in_buf[574]*(-14)+in_buf[575]*(2)+in_buf[576]*(-20)+in_buf[577]*(-15)+in_buf[578]*(-15)+in_buf[579]*(-9)+in_buf[580]*(5)+in_buf[581]*(9)+in_buf[582]*(13)+in_buf[583]*(8)+in_buf[584]*(-7)+in_buf[585]*(-6)+in_buf[586]*(-50)+in_buf[587]*(0)+in_buf[588]*(-2)+in_buf[589]*(-3)+in_buf[590]*(-7)+in_buf[591]*(-27)+in_buf[592]*(-22)+in_buf[593]*(-16)+in_buf[594]*(-13)+in_buf[595]*(0)+in_buf[596]*(6)+in_buf[597]*(3)+in_buf[598]*(-16)+in_buf[599]*(0)+in_buf[600]*(-12)+in_buf[601]*(-8)+in_buf[602]*(-7)+in_buf[603]*(6)+in_buf[604]*(-13)+in_buf[605]*(-12)+in_buf[606]*(-14)+in_buf[607]*(-3)+in_buf[608]*(5)+in_buf[609]*(12)+in_buf[610]*(9)+in_buf[611]*(13)+in_buf[612]*(1)+in_buf[613]*(3)+in_buf[614]*(-23)+in_buf[615]*(-2)+in_buf[616]*(-5)+in_buf[617]*(2)+in_buf[618]*(-6)+in_buf[619]*(3)+in_buf[620]*(7)+in_buf[621]*(-29)+in_buf[622]*(-19)+in_buf[623]*(1)+in_buf[624]*(-5)+in_buf[625]*(-6)+in_buf[626]*(-6)+in_buf[627]*(2)+in_buf[628]*(0)+in_buf[629]*(-4)+in_buf[630]*(2)+in_buf[631]*(3)+in_buf[632]*(-4)+in_buf[633]*(-3)+in_buf[634]*(1)+in_buf[635]*(8)+in_buf[636]*(8)+in_buf[637]*(9)+in_buf[638]*(4)+in_buf[639]*(27)+in_buf[640]*(4)+in_buf[641]*(4)+in_buf[642]*(17)+in_buf[643]*(1)+in_buf[644]*(-3)+in_buf[645]*(-3)+in_buf[646]*(9)+in_buf[647]*(19)+in_buf[648]*(32)+in_buf[649]*(-5)+in_buf[650]*(-9)+in_buf[651]*(-15)+in_buf[652]*(4)+in_buf[653]*(-5)+in_buf[654]*(9)+in_buf[655]*(6)+in_buf[656]*(4)+in_buf[657]*(10)+in_buf[658]*(11)+in_buf[659]*(8)+in_buf[660]*(8)+in_buf[661]*(1)+in_buf[662]*(17)+in_buf[663]*(14)+in_buf[664]*(5)+in_buf[665]*(4)+in_buf[666]*(9)+in_buf[667]*(14)+in_buf[668]*(3)+in_buf[669]*(8)+in_buf[670]*(18)+in_buf[671]*(-2)+in_buf[672]*(2)+in_buf[673]*(1)+in_buf[674]*(-17)+in_buf[675]*(-5)+in_buf[676]*(-8)+in_buf[677]*(0)+in_buf[678]*(-4)+in_buf[679]*(12)+in_buf[680]*(13)+in_buf[681]*(6)+in_buf[682]*(19)+in_buf[683]*(38)+in_buf[684]*(21)+in_buf[685]*(21)+in_buf[686]*(21)+in_buf[687]*(17)+in_buf[688]*(23)+in_buf[689]*(-5)+in_buf[690]*(7)+in_buf[691]*(30)+in_buf[692]*(19)+in_buf[693]*(13)+in_buf[694]*(0)+in_buf[695]*(-15)+in_buf[696]*(-29)+in_buf[697]*(-14)+in_buf[698]*(-14)+in_buf[699]*(0)+in_buf[700]*(3)+in_buf[701]*(4)+in_buf[702]*(21)+in_buf[703]*(1)+in_buf[704]*(-45)+in_buf[705]*(-40)+in_buf[706]*(0)+in_buf[707]*(15)+in_buf[708]*(-16)+in_buf[709]*(4)+in_buf[710]*(35)+in_buf[711]*(21)+in_buf[712]*(13)+in_buf[713]*(32)+in_buf[714]*(20)+in_buf[715]*(32)+in_buf[716]*(27)+in_buf[717]*(32)+in_buf[718]*(37)+in_buf[719]*(32)+in_buf[720]*(19)+in_buf[721]*(36)+in_buf[722]*(43)+in_buf[723]*(42)+in_buf[724]*(25)+in_buf[725]*(2)+in_buf[726]*(-12)+in_buf[727]*(-2)+in_buf[728]*(3)+in_buf[729]*(4)+in_buf[730]*(0)+in_buf[731]*(-16)+in_buf[732]*(-42)+in_buf[733]*(-22)+in_buf[734]*(-39)+in_buf[735]*(-37)+in_buf[736]*(10)+in_buf[737]*(-5)+in_buf[738]*(-1)+in_buf[739]*(13)+in_buf[740]*(9)+in_buf[741]*(-9)+in_buf[742]*(-18)+in_buf[743]*(-2)+in_buf[744]*(19)+in_buf[745]*(10)+in_buf[746]*(-13)+in_buf[747]*(-36)+in_buf[748]*(-47)+in_buf[749]*(-23)+in_buf[750]*(2)+in_buf[751]*(7)+in_buf[752]*(-16)+in_buf[753]*(0)+in_buf[754]*(4)+in_buf[755]*(-1)+in_buf[756]*(4)+in_buf[757]*(-3)+in_buf[758]*(1)+in_buf[759]*(0)+in_buf[760]*(-18)+in_buf[761]*(-27)+in_buf[762]*(-19)+in_buf[763]*(-5)+in_buf[764]*(-11)+in_buf[765]*(-26)+in_buf[766]*(-43)+in_buf[767]*(-20)+in_buf[768]*(-14)+in_buf[769]*(-40)+in_buf[770]*(-60)+in_buf[771]*(-6)+in_buf[772]*(-21)+in_buf[773]*(-42)+in_buf[774]*(-26)+in_buf[775]*(-20)+in_buf[776]*(-2)+in_buf[777]*(-16)+in_buf[778]*(8)+in_buf[779]*(-1)+in_buf[780]*(-2)+in_buf[781]*(0)+in_buf[782]*(-3)+in_buf[783]*(4);
assign in_buf_weight033=in_buf[0]*(1)+in_buf[1]*(2)+in_buf[2]*(-2)+in_buf[3]*(1)+in_buf[4]*(-2)+in_buf[5]*(1)+in_buf[6]*(0)+in_buf[7]*(4)+in_buf[8]*(2)+in_buf[9]*(-2)+in_buf[10]*(4)+in_buf[11]*(2)+in_buf[12]*(-10)+in_buf[13]*(0)+in_buf[14]*(29)+in_buf[15]*(15)+in_buf[16]*(3)+in_buf[17]*(0)+in_buf[18]*(2)+in_buf[19]*(3)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(4)+in_buf[23]*(1)+in_buf[24]*(0)+in_buf[25]*(1)+in_buf[26]*(-3)+in_buf[27]*(-2)+in_buf[28]*(-1)+in_buf[29]*(0)+in_buf[30]*(3)+in_buf[31]*(-2)+in_buf[32]*(-2)+in_buf[33]*(4)+in_buf[34]*(0)+in_buf[35]*(-7)+in_buf[36]*(2)+in_buf[37]*(6)+in_buf[38]*(9)+in_buf[39]*(24)+in_buf[40]*(6)+in_buf[41]*(13)+in_buf[42]*(-17)+in_buf[43]*(5)+in_buf[44]*(34)+in_buf[45]*(26)+in_buf[46]*(-28)+in_buf[47]*(-27)+in_buf[48]*(-37)+in_buf[49]*(-23)+in_buf[50]*(-24)+in_buf[51]*(-17)+in_buf[52]*(0)+in_buf[53]*(3)+in_buf[54]*(-1)+in_buf[55]*(-3)+in_buf[56]*(-3)+in_buf[57]*(0)+in_buf[58]*(-2)+in_buf[59]*(31)+in_buf[60]*(30)+in_buf[61]*(-3)+in_buf[62]*(-4)+in_buf[63]*(3)+in_buf[64]*(11)+in_buf[65]*(33)+in_buf[66]*(31)+in_buf[67]*(13)+in_buf[68]*(-28)+in_buf[69]*(-44)+in_buf[70]*(-31)+in_buf[71]*(-34)+in_buf[72]*(-17)+in_buf[73]*(17)+in_buf[74]*(20)+in_buf[75]*(18)+in_buf[76]*(7)+in_buf[77]*(-2)+in_buf[78]*(-24)+in_buf[79]*(2)+in_buf[80]*(12)+in_buf[81]*(10)+in_buf[82]*(0)+in_buf[83]*(0)+in_buf[84]*(-3)+in_buf[85]*(-1)+in_buf[86]*(-12)+in_buf[87]*(23)+in_buf[88]*(26)+in_buf[89]*(16)+in_buf[90]*(-3)+in_buf[91]*(-42)+in_buf[92]*(-16)+in_buf[93]*(8)+in_buf[94]*(0)+in_buf[95]*(33)+in_buf[96]*(-1)+in_buf[97]*(-37)+in_buf[98]*(-17)+in_buf[99]*(-18)+in_buf[100]*(-21)+in_buf[101]*(11)+in_buf[102]*(-4)+in_buf[103]*(-6)+in_buf[104]*(18)+in_buf[105]*(21)+in_buf[106]*(11)+in_buf[107]*(-6)+in_buf[108]*(26)+in_buf[109]*(44)+in_buf[110]*(38)+in_buf[111]*(-3)+in_buf[112]*(-1)+in_buf[113]*(-4)+in_buf[114]*(-22)+in_buf[115]*(-9)+in_buf[116]*(-22)+in_buf[117]*(-8)+in_buf[118]*(-26)+in_buf[119]*(-45)+in_buf[120]*(-52)+in_buf[121]*(-44)+in_buf[122]*(-49)+in_buf[123]*(-20)+in_buf[124]*(-33)+in_buf[125]*(-48)+in_buf[126]*(-38)+in_buf[127]*(-21)+in_buf[128]*(-7)+in_buf[129]*(7)+in_buf[130]*(16)+in_buf[131]*(1)+in_buf[132]*(0)+in_buf[133]*(8)+in_buf[134]*(-4)+in_buf[135]*(20)+in_buf[136]*(41)+in_buf[137]*(27)+in_buf[138]*(-4)+in_buf[139]*(8)+in_buf[140]*(-3)+in_buf[141]*(4)+in_buf[142]*(-29)+in_buf[143]*(-15)+in_buf[144]*(-46)+in_buf[145]*(-28)+in_buf[146]*(-50)+in_buf[147]*(-68)+in_buf[148]*(-31)+in_buf[149]*(-26)+in_buf[150]*(-55)+in_buf[151]*(-23)+in_buf[152]*(-29)+in_buf[153]*(-19)+in_buf[154]*(-13)+in_buf[155]*(-19)+in_buf[156]*(-16)+in_buf[157]*(-10)+in_buf[158]*(-6)+in_buf[159]*(-14)+in_buf[160]*(-13)+in_buf[161]*(-7)+in_buf[162]*(-8)+in_buf[163]*(-3)+in_buf[164]*(7)+in_buf[165]*(16)+in_buf[166]*(-10)+in_buf[167]*(15)+in_buf[168]*(0)+in_buf[169]*(-24)+in_buf[170]*(16)+in_buf[171]*(-4)+in_buf[172]*(18)+in_buf[173]*(6)+in_buf[174]*(-12)+in_buf[175]*(-6)+in_buf[176]*(8)+in_buf[177]*(0)+in_buf[178]*(-11)+in_buf[179]*(3)+in_buf[180]*(-13)+in_buf[181]*(-3)+in_buf[182]*(-6)+in_buf[183]*(-16)+in_buf[184]*(-11)+in_buf[185]*(-6)+in_buf[186]*(-9)+in_buf[187]*(-4)+in_buf[188]*(-14)+in_buf[189]*(-4)+in_buf[190]*(0)+in_buf[191]*(-11)+in_buf[192]*(2)+in_buf[193]*(-2)+in_buf[194]*(0)+in_buf[195]*(-10)+in_buf[196]*(1)+in_buf[197]*(-9)+in_buf[198]*(29)+in_buf[199]*(22)+in_buf[200]*(-3)+in_buf[201]*(-3)+in_buf[202]*(6)+in_buf[203]*(-6)+in_buf[204]*(4)+in_buf[205]*(7)+in_buf[206]*(-5)+in_buf[207]*(3)+in_buf[208]*(-7)+in_buf[209]*(4)+in_buf[210]*(4)+in_buf[211]*(-2)+in_buf[212]*(4)+in_buf[213]*(3)+in_buf[214]*(0)+in_buf[215]*(-1)+in_buf[216]*(4)+in_buf[217]*(2)+in_buf[218]*(-11)+in_buf[219]*(-7)+in_buf[220]*(7)+in_buf[221]*(14)+in_buf[222]*(9)+in_buf[223]*(3)+in_buf[224]*(11)+in_buf[225]*(38)+in_buf[226]*(22)+in_buf[227]*(-19)+in_buf[228]*(-25)+in_buf[229]*(-3)+in_buf[230]*(3)+in_buf[231]*(-7)+in_buf[232]*(0)+in_buf[233]*(-5)+in_buf[234]*(-6)+in_buf[235]*(-5)+in_buf[236]*(-1)+in_buf[237]*(3)+in_buf[238]*(2)+in_buf[239]*(18)+in_buf[240]*(12)+in_buf[241]*(5)+in_buf[242]*(0)+in_buf[243]*(1)+in_buf[244]*(13)+in_buf[245]*(0)+in_buf[246]*(-17)+in_buf[247]*(6)+in_buf[248]*(28)+in_buf[249]*(21)+in_buf[250]*(-15)+in_buf[251]*(0)+in_buf[252]*(10)+in_buf[253]*(33)+in_buf[254]*(-2)+in_buf[255]*(1)+in_buf[256]*(-20)+in_buf[257]*(-4)+in_buf[258]*(-6)+in_buf[259]*(-6)+in_buf[260]*(-16)+in_buf[261]*(-26)+in_buf[262]*(0)+in_buf[263]*(10)+in_buf[264]*(30)+in_buf[265]*(25)+in_buf[266]*(20)+in_buf[267]*(14)+in_buf[268]*(10)+in_buf[269]*(12)+in_buf[270]*(10)+in_buf[271]*(11)+in_buf[272]*(9)+in_buf[273]*(-11)+in_buf[274]*(-17)+in_buf[275]*(-6)+in_buf[276]*(34)+in_buf[277]*(3)+in_buf[278]*(6)+in_buf[279]*(22)+in_buf[280]*(13)+in_buf[281]*(16)+in_buf[282]*(35)+in_buf[283]*(8)+in_buf[284]*(-21)+in_buf[285]*(3)+in_buf[286]*(12)+in_buf[287]*(0)+in_buf[288]*(-16)+in_buf[289]*(-4)+in_buf[290]*(14)+in_buf[291]*(25)+in_buf[292]*(36)+in_buf[293]*(31)+in_buf[294]*(27)+in_buf[295]*(20)+in_buf[296]*(16)+in_buf[297]*(14)+in_buf[298]*(16)+in_buf[299]*(19)+in_buf[300]*(19)+in_buf[301]*(1)+in_buf[302]*(-16)+in_buf[303]*(-8)+in_buf[304]*(41)+in_buf[305]*(45)+in_buf[306]*(32)+in_buf[307]*(-1)+in_buf[308]*(12)+in_buf[309]*(46)+in_buf[310]*(24)+in_buf[311]*(-5)+in_buf[312]*(-18)+in_buf[313]*(-24)+in_buf[314]*(6)+in_buf[315]*(-14)+in_buf[316]*(-14)+in_buf[317]*(-5)+in_buf[318]*(5)+in_buf[319]*(19)+in_buf[320]*(26)+in_buf[321]*(16)+in_buf[322]*(2)+in_buf[323]*(4)+in_buf[324]*(-7)+in_buf[325]*(0)+in_buf[326]*(12)+in_buf[327]*(19)+in_buf[328]*(5)+in_buf[329]*(-13)+in_buf[330]*(-11)+in_buf[331]*(-6)+in_buf[332]*(8)+in_buf[333]*(31)+in_buf[334]*(-3)+in_buf[335]*(-2)+in_buf[336]*(21)+in_buf[337]*(13)+in_buf[338]*(31)+in_buf[339]*(6)+in_buf[340]*(-10)+in_buf[341]*(-13)+in_buf[342]*(-7)+in_buf[343]*(-6)+in_buf[344]*(9)+in_buf[345]*(7)+in_buf[346]*(5)+in_buf[347]*(16)+in_buf[348]*(26)+in_buf[349]*(15)+in_buf[350]*(10)+in_buf[351]*(-1)+in_buf[352]*(-13)+in_buf[353]*(-5)+in_buf[354]*(13)+in_buf[355]*(2)+in_buf[356]*(-11)+in_buf[357]*(-30)+in_buf[358]*(-17)+in_buf[359]*(-44)+in_buf[360]*(-40)+in_buf[361]*(12)+in_buf[362]*(7)+in_buf[363]*(11)+in_buf[364]*(-5)+in_buf[365]*(1)+in_buf[366]*(44)+in_buf[367]*(36)+in_buf[368]*(13)+in_buf[369]*(13)+in_buf[370]*(16)+in_buf[371]*(18)+in_buf[372]*(3)+in_buf[373]*(-1)+in_buf[374]*(18)+in_buf[375]*(21)+in_buf[376]*(26)+in_buf[377]*(12)+in_buf[378]*(1)+in_buf[379]*(-4)+in_buf[380]*(-7)+in_buf[381]*(-3)+in_buf[382]*(-1)+in_buf[383]*(-7)+in_buf[384]*(-20)+in_buf[385]*(-19)+in_buf[386]*(-23)+in_buf[387]*(-29)+in_buf[388]*(-15)+in_buf[389]*(-13)+in_buf[390]*(3)+in_buf[391]*(19)+in_buf[392]*(16)+in_buf[393]*(4)+in_buf[394]*(20)+in_buf[395]*(57)+in_buf[396]*(39)+in_buf[397]*(27)+in_buf[398]*(26)+in_buf[399]*(29)+in_buf[400]*(0)+in_buf[401]*(-4)+in_buf[402]*(5)+in_buf[403]*(5)+in_buf[404]*(10)+in_buf[405]*(-1)+in_buf[406]*(-4)+in_buf[407]*(-4)+in_buf[408]*(0)+in_buf[409]*(18)+in_buf[410]*(11)+in_buf[411]*(-12)+in_buf[412]*(-10)+in_buf[413]*(-21)+in_buf[414]*(-6)+in_buf[415]*(7)+in_buf[416]*(20)+in_buf[417]*(-6)+in_buf[418]*(19)+in_buf[419]*(23)+in_buf[420]*(19)+in_buf[421]*(-4)+in_buf[422]*(-14)+in_buf[423]*(60)+in_buf[424]*(45)+in_buf[425]*(32)+in_buf[426]*(26)+in_buf[427]*(8)+in_buf[428]*(-23)+in_buf[429]*(-9)+in_buf[430]*(8)+in_buf[431]*(11)+in_buf[432]*(19)+in_buf[433]*(-17)+in_buf[434]*(-7)+in_buf[435]*(7)+in_buf[436]*(15)+in_buf[437]*(33)+in_buf[438]*(26)+in_buf[439]*(-8)+in_buf[440]*(-9)+in_buf[441]*(-1)+in_buf[442]*(9)+in_buf[443]*(28)+in_buf[444]*(38)+in_buf[445]*(2)+in_buf[446]*(9)+in_buf[447]*(28)+in_buf[448]*(3)+in_buf[449]*(-24)+in_buf[450]*(-21)+in_buf[451]*(23)+in_buf[452]*(23)+in_buf[453]*(22)+in_buf[454]*(8)+in_buf[455]*(7)+in_buf[456]*(-4)+in_buf[457]*(-17)+in_buf[458]*(-6)+in_buf[459]*(2)+in_buf[460]*(11)+in_buf[461]*(-2)+in_buf[462]*(-6)+in_buf[463]*(17)+in_buf[464]*(22)+in_buf[465]*(43)+in_buf[466]*(22)+in_buf[467]*(14)+in_buf[468]*(5)+in_buf[469]*(17)+in_buf[470]*(16)+in_buf[471]*(16)+in_buf[472]*(-10)+in_buf[473]*(6)+in_buf[474]*(36)+in_buf[475]*(30)+in_buf[476]*(2)+in_buf[477]*(-12)+in_buf[478]*(-8)+in_buf[479]*(-4)+in_buf[480]*(9)+in_buf[481]*(31)+in_buf[482]*(25)+in_buf[483]*(1)+in_buf[484]*(5)+in_buf[485]*(12)+in_buf[486]*(-4)+in_buf[487]*(-6)+in_buf[488]*(-9)+in_buf[489]*(-9)+in_buf[490]*(5)+in_buf[491]*(21)+in_buf[492]*(26)+in_buf[493]*(31)+in_buf[494]*(11)+in_buf[495]*(0)+in_buf[496]*(15)+in_buf[497]*(12)+in_buf[498]*(-4)+in_buf[499]*(-19)+in_buf[500]*(-30)+in_buf[501]*(1)+in_buf[502]*(12)+in_buf[503]*(27)+in_buf[504]*(10)+in_buf[505]*(-13)+in_buf[506]*(-6)+in_buf[507]*(-15)+in_buf[508]*(5)+in_buf[509]*(32)+in_buf[510]*(23)+in_buf[511]*(8)+in_buf[512]*(16)+in_buf[513]*(-4)+in_buf[514]*(-7)+in_buf[515]*(-4)+in_buf[516]*(-17)+in_buf[517]*(-4)+in_buf[518]*(6)+in_buf[519]*(3)+in_buf[520]*(20)+in_buf[521]*(18)+in_buf[522]*(6)+in_buf[523]*(6)+in_buf[524]*(11)+in_buf[525]*(-7)+in_buf[526]*(-9)+in_buf[527]*(-13)+in_buf[528]*(-12)+in_buf[529]*(-10)+in_buf[530]*(0)+in_buf[531]*(5)+in_buf[532]*(-8)+in_buf[533]*(18)+in_buf[534]*(1)+in_buf[535]*(0)+in_buf[536]*(-3)+in_buf[537]*(5)+in_buf[538]*(9)+in_buf[539]*(2)+in_buf[540]*(6)+in_buf[541]*(-3)+in_buf[542]*(5)+in_buf[543]*(1)+in_buf[544]*(-1)+in_buf[545]*(-2)+in_buf[546]*(7)+in_buf[547]*(0)+in_buf[548]*(4)+in_buf[549]*(7)+in_buf[550]*(7)+in_buf[551]*(3)+in_buf[552]*(10)+in_buf[553]*(-9)+in_buf[554]*(-8)+in_buf[555]*(1)+in_buf[556]*(-12)+in_buf[557]*(-16)+in_buf[558]*(31)+in_buf[559]*(-12)+in_buf[560]*(-1)+in_buf[561]*(26)+in_buf[562]*(8)+in_buf[563]*(15)+in_buf[564]*(2)+in_buf[565]*(0)+in_buf[566]*(0)+in_buf[567]*(-12)+in_buf[568]*(9)+in_buf[569]*(13)+in_buf[570]*(12)+in_buf[571]*(10)+in_buf[572]*(2)+in_buf[573]*(-3)+in_buf[574]*(-10)+in_buf[575]*(-22)+in_buf[576]*(-23)+in_buf[577]*(-4)+in_buf[578]*(-4)+in_buf[579]*(-12)+in_buf[580]*(-14)+in_buf[581]*(-23)+in_buf[582]*(-26)+in_buf[583]*(-18)+in_buf[584]*(8)+in_buf[585]*(17)+in_buf[586]*(20)+in_buf[587]*(0)+in_buf[588]*(-1)+in_buf[589]*(-10)+in_buf[590]*(4)+in_buf[591]*(3)+in_buf[592]*(2)+in_buf[593]*(4)+in_buf[594]*(-7)+in_buf[595]*(-3)+in_buf[596]*(-1)+in_buf[597]*(2)+in_buf[598]*(-5)+in_buf[599]*(-7)+in_buf[600]*(-4)+in_buf[601]*(-9)+in_buf[602]*(-24)+in_buf[603]*(-31)+in_buf[604]*(-18)+in_buf[605]*(-3)+in_buf[606]*(-2)+in_buf[607]*(-18)+in_buf[608]*(-35)+in_buf[609]*(-29)+in_buf[610]*(-34)+in_buf[611]*(-29)+in_buf[612]*(2)+in_buf[613]*(26)+in_buf[614]*(39)+in_buf[615]*(4)+in_buf[616]*(2)+in_buf[617]*(-13)+in_buf[618]*(-14)+in_buf[619]*(23)+in_buf[620]*(-10)+in_buf[621]*(-23)+in_buf[622]*(-10)+in_buf[623]*(7)+in_buf[624]*(5)+in_buf[625]*(2)+in_buf[626]*(0)+in_buf[627]*(-14)+in_buf[628]*(-1)+in_buf[629]*(-23)+in_buf[630]*(-28)+in_buf[631]*(-22)+in_buf[632]*(-3)+in_buf[633]*(0)+in_buf[634]*(-10)+in_buf[635]*(-29)+in_buf[636]*(-36)+in_buf[637]*(-41)+in_buf[638]*(-31)+in_buf[639]*(-4)+in_buf[640]*(39)+in_buf[641]*(24)+in_buf[642]*(8)+in_buf[643]*(1)+in_buf[644]*(-2)+in_buf[645]*(5)+in_buf[646]*(-36)+in_buf[647]*(33)+in_buf[648]*(2)+in_buf[649]*(-17)+in_buf[650]*(15)+in_buf[651]*(16)+in_buf[652]*(4)+in_buf[653]*(-6)+in_buf[654]*(0)+in_buf[655]*(-13)+in_buf[656]*(-24)+in_buf[657]*(-41)+in_buf[658]*(-34)+in_buf[659]*(-31)+in_buf[660]*(-5)+in_buf[661]*(-3)+in_buf[662]*(-15)+in_buf[663]*(-28)+in_buf[664]*(-47)+in_buf[665]*(-36)+in_buf[666]*(7)+in_buf[667]*(12)+in_buf[668]*(55)+in_buf[669]*(20)+in_buf[670]*(-1)+in_buf[671]*(0)+in_buf[672]*(2)+in_buf[673]*(4)+in_buf[674]*(-16)+in_buf[675]*(3)+in_buf[676]*(9)+in_buf[677]*(-5)+in_buf[678]*(-1)+in_buf[679]*(6)+in_buf[680]*(1)+in_buf[681]*(1)+in_buf[682]*(-17)+in_buf[683]*(-21)+in_buf[684]*(-28)+in_buf[685]*(-19)+in_buf[686]*(-26)+in_buf[687]*(-29)+in_buf[688]*(-6)+in_buf[689]*(15)+in_buf[690]*(4)+in_buf[691]*(-18)+in_buf[692]*(-15)+in_buf[693]*(11)+in_buf[694]*(45)+in_buf[695]*(40)+in_buf[696]*(39)+in_buf[697]*(1)+in_buf[698]*(10)+in_buf[699]*(0)+in_buf[700]*(-1)+in_buf[701]*(3)+in_buf[702]*(9)+in_buf[703]*(15)+in_buf[704]*(1)+in_buf[705]*(-1)+in_buf[706]*(-15)+in_buf[707]*(-1)+in_buf[708]*(-20)+in_buf[709]*(-21)+in_buf[710]*(-22)+in_buf[711]*(10)+in_buf[712]*(-6)+in_buf[713]*(14)+in_buf[714]*(-7)+in_buf[715]*(4)+in_buf[716]*(20)+in_buf[717]*(27)+in_buf[718]*(12)+in_buf[719]*(12)+in_buf[720]*(26)+in_buf[721]*(70)+in_buf[722]*(81)+in_buf[723]*(58)+in_buf[724]*(44)+in_buf[725]*(25)+in_buf[726]*(8)+in_buf[727]*(2)+in_buf[728]*(0)+in_buf[729]*(-1)+in_buf[730]*(3)+in_buf[731]*(10)+in_buf[732]*(-5)+in_buf[733]*(-19)+in_buf[734]*(-21)+in_buf[735]*(-9)+in_buf[736]*(0)+in_buf[737]*(-4)+in_buf[738]*(-12)+in_buf[739]*(21)+in_buf[740]*(27)+in_buf[741]*(43)+in_buf[742]*(37)+in_buf[743]*(38)+in_buf[744]*(24)+in_buf[745]*(-1)+in_buf[746]*(1)+in_buf[747]*(51)+in_buf[748]*(35)+in_buf[749]*(33)+in_buf[750]*(43)+in_buf[751]*(-22)+in_buf[752]*(-32)+in_buf[753]*(14)+in_buf[754]*(2)+in_buf[755]*(1)+in_buf[756]*(4)+in_buf[757]*(2)+in_buf[758]*(0)+in_buf[759]*(1)+in_buf[760]*(16)+in_buf[761]*(18)+in_buf[762]*(10)+in_buf[763]*(7)+in_buf[764]*(11)+in_buf[765]*(22)+in_buf[766]*(27)+in_buf[767]*(24)+in_buf[768]*(21)+in_buf[769]*(38)+in_buf[770]*(33)+in_buf[771]*(8)+in_buf[772]*(16)+in_buf[773]*(34)+in_buf[774]*(33)+in_buf[775]*(28)+in_buf[776]*(41)+in_buf[777]*(36)+in_buf[778]*(33)+in_buf[779]*(9)+in_buf[780]*(-3)+in_buf[781]*(1)+in_buf[782]*(-2)+in_buf[783]*(-3);
assign in_buf_weight034=in_buf[0]*(0)+in_buf[1]*(4)+in_buf[2]*(-1)+in_buf[3]*(2)+in_buf[4]*(0)+in_buf[5]*(0)+in_buf[6]*(2)+in_buf[7]*(3)+in_buf[8]*(0)+in_buf[9]*(-2)+in_buf[10]*(-1)+in_buf[11]*(-1)+in_buf[12]*(-4)+in_buf[13]*(-9)+in_buf[14]*(0)+in_buf[15]*(2)+in_buf[16]*(2)+in_buf[17]*(0)+in_buf[18]*(-1)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(3)+in_buf[22]*(0)+in_buf[23]*(-3)+in_buf[24]*(4)+in_buf[25]*(2)+in_buf[26]*(-1)+in_buf[27]*(1)+in_buf[28]*(0)+in_buf[29]*(-1)+in_buf[30]*(-2)+in_buf[31]*(1)+in_buf[32]*(0)+in_buf[33]*(-2)+in_buf[34]*(1)+in_buf[35]*(0)+in_buf[36]*(-5)+in_buf[37]*(1)+in_buf[38]*(-10)+in_buf[39]*(6)+in_buf[40]*(8)+in_buf[41]*(13)+in_buf[42]*(44)+in_buf[43]*(36)+in_buf[44]*(31)+in_buf[45]*(10)+in_buf[46]*(-24)+in_buf[47]*(-14)+in_buf[48]*(-15)+in_buf[49]*(-30)+in_buf[50]*(-24)+in_buf[51]*(-13)+in_buf[52]*(0)+in_buf[53]*(-1)+in_buf[54]*(2)+in_buf[55]*(-3)+in_buf[56]*(1)+in_buf[57]*(0)+in_buf[58]*(-6)+in_buf[59]*(30)+in_buf[60]*(28)+in_buf[61]*(-3)+in_buf[62]*(-2)+in_buf[63]*(-4)+in_buf[64]*(-7)+in_buf[65]*(-11)+in_buf[66]*(-27)+in_buf[67]*(-37)+in_buf[68]*(-17)+in_buf[69]*(16)+in_buf[70]*(2)+in_buf[71]*(-27)+in_buf[72]*(-16)+in_buf[73]*(-25)+in_buf[74]*(-36)+in_buf[75]*(-30)+in_buf[76]*(-45)+in_buf[77]*(-40)+in_buf[78]*(-33)+in_buf[79]*(-23)+in_buf[80]*(0)+in_buf[81]*(2)+in_buf[82]*(3)+in_buf[83]*(0)+in_buf[84]*(3)+in_buf[85]*(0)+in_buf[86]*(7)+in_buf[87]*(26)+in_buf[88]*(12)+in_buf[89]*(-24)+in_buf[90]*(-23)+in_buf[91]*(-14)+in_buf[92]*(-14)+in_buf[93]*(-4)+in_buf[94]*(-26)+in_buf[95]*(-35)+in_buf[96]*(-34)+in_buf[97]*(-46)+in_buf[98]*(-52)+in_buf[99]*(-32)+in_buf[100]*(-25)+in_buf[101]*(-25)+in_buf[102]*(-38)+in_buf[103]*(-45)+in_buf[104]*(-30)+in_buf[105]*(-13)+in_buf[106]*(-21)+in_buf[107]*(-21)+in_buf[108]*(0)+in_buf[109]*(8)+in_buf[110]*(6)+in_buf[111]*(-3)+in_buf[112]*(0)+in_buf[113]*(3)+in_buf[114]*(6)+in_buf[115]*(14)+in_buf[116]*(4)+in_buf[117]*(-24)+in_buf[118]*(-36)+in_buf[119]*(-33)+in_buf[120]*(-42)+in_buf[121]*(-16)+in_buf[122]*(-22)+in_buf[123]*(-11)+in_buf[124]*(-15)+in_buf[125]*(-29)+in_buf[126]*(-11)+in_buf[127]*(-2)+in_buf[128]*(-19)+in_buf[129]*(-8)+in_buf[130]*(-23)+in_buf[131]*(-32)+in_buf[132]*(-10)+in_buf[133]*(7)+in_buf[134]*(-29)+in_buf[135]*(-33)+in_buf[136]*(-10)+in_buf[137]*(5)+in_buf[138]*(2)+in_buf[139]*(-15)+in_buf[140]*(-3)+in_buf[141]*(0)+in_buf[142]*(0)+in_buf[143]*(-9)+in_buf[144]*(-18)+in_buf[145]*(-22)+in_buf[146]*(-34)+in_buf[147]*(-27)+in_buf[148]*(-18)+in_buf[149]*(-21)+in_buf[150]*(-10)+in_buf[151]*(1)+in_buf[152]*(-2)+in_buf[153]*(-5)+in_buf[154]*(-16)+in_buf[155]*(-9)+in_buf[156]*(-29)+in_buf[157]*(-31)+in_buf[158]*(-39)+in_buf[159]*(-31)+in_buf[160]*(-17)+in_buf[161]*(-3)+in_buf[162]*(-35)+in_buf[163]*(-43)+in_buf[164]*(-28)+in_buf[165]*(-16)+in_buf[166]*(-8)+in_buf[167]*(-13)+in_buf[168]*(3)+in_buf[169]*(-13)+in_buf[170]*(-2)+in_buf[171]*(4)+in_buf[172]*(-13)+in_buf[173]*(-30)+in_buf[174]*(-23)+in_buf[175]*(-18)+in_buf[176]*(-22)+in_buf[177]*(-9)+in_buf[178]*(4)+in_buf[179]*(0)+in_buf[180]*(0)+in_buf[181]*(13)+in_buf[182]*(13)+in_buf[183]*(-4)+in_buf[184]*(-9)+in_buf[185]*(-9)+in_buf[186]*(-16)+in_buf[187]*(-26)+in_buf[188]*(-12)+in_buf[189]*(-1)+in_buf[190]*(-8)+in_buf[191]*(-21)+in_buf[192]*(-23)+in_buf[193]*(-16)+in_buf[194]*(-10)+in_buf[195]*(-10)+in_buf[196]*(5)+in_buf[197]*(-28)+in_buf[198]*(0)+in_buf[199]*(11)+in_buf[200]*(-17)+in_buf[201]*(-39)+in_buf[202]*(-26)+in_buf[203]*(-24)+in_buf[204]*(-11)+in_buf[205]*(-3)+in_buf[206]*(17)+in_buf[207]*(6)+in_buf[208]*(3)+in_buf[209]*(1)+in_buf[210]*(-3)+in_buf[211]*(10)+in_buf[212]*(16)+in_buf[213]*(-2)+in_buf[214]*(-2)+in_buf[215]*(-8)+in_buf[216]*(-11)+in_buf[217]*(-4)+in_buf[218]*(-1)+in_buf[219]*(-1)+in_buf[220]*(-7)+in_buf[221]*(0)+in_buf[222]*(-14)+in_buf[223]*(-2)+in_buf[224]*(-30)+in_buf[225]*(16)+in_buf[226]*(-25)+in_buf[227]*(-16)+in_buf[228]*(-18)+in_buf[229]*(-23)+in_buf[230]*(-5)+in_buf[231]*(-6)+in_buf[232]*(3)+in_buf[233]*(-6)+in_buf[234]*(7)+in_buf[235]*(1)+in_buf[236]*(0)+in_buf[237]*(2)+in_buf[238]*(10)+in_buf[239]*(19)+in_buf[240]*(33)+in_buf[241]*(18)+in_buf[242]*(17)+in_buf[243]*(12)+in_buf[244]*(0)+in_buf[245]*(2)+in_buf[246]*(2)+in_buf[247]*(2)+in_buf[248]*(33)+in_buf[249]*(10)+in_buf[250]*(-13)+in_buf[251]*(27)+in_buf[252]*(6)+in_buf[253]*(26)+in_buf[254]*(-10)+in_buf[255]*(1)+in_buf[256]*(-12)+in_buf[257]*(-16)+in_buf[258]*(-1)+in_buf[259]*(-10)+in_buf[260]*(-11)+in_buf[261]*(2)+in_buf[262]*(23)+in_buf[263]*(9)+in_buf[264]*(1)+in_buf[265]*(15)+in_buf[266]*(22)+in_buf[267]*(24)+in_buf[268]*(22)+in_buf[269]*(24)+in_buf[270]*(23)+in_buf[271]*(5)+in_buf[272]*(-5)+in_buf[273]*(-3)+in_buf[274]*(4)+in_buf[275]*(-4)+in_buf[276]*(19)+in_buf[277]*(30)+in_buf[278]*(19)+in_buf[279]*(32)+in_buf[280]*(3)+in_buf[281]*(9)+in_buf[282]*(14)+in_buf[283]*(4)+in_buf[284]*(-13)+in_buf[285]*(-16)+in_buf[286]*(-4)+in_buf[287]*(-8)+in_buf[288]*(-7)+in_buf[289]*(3)+in_buf[290]*(9)+in_buf[291]*(1)+in_buf[292]*(0)+in_buf[293]*(9)+in_buf[294]*(29)+in_buf[295]*(38)+in_buf[296]*(24)+in_buf[297]*(10)+in_buf[298]*(12)+in_buf[299]*(5)+in_buf[300]*(1)+in_buf[301]*(2)+in_buf[302]*(19)+in_buf[303]*(19)+in_buf[304]*(28)+in_buf[305]*(59)+in_buf[306]*(39)+in_buf[307]*(22)+in_buf[308]*(5)+in_buf[309]*(-27)+in_buf[310]*(38)+in_buf[311]*(22)+in_buf[312]*(-3)+in_buf[313]*(-11)+in_buf[314]*(2)+in_buf[315]*(0)+in_buf[316]*(4)+in_buf[317]*(-3)+in_buf[318]*(-2)+in_buf[319]*(0)+in_buf[320]*(-1)+in_buf[321]*(23)+in_buf[322]*(52)+in_buf[323]*(37)+in_buf[324]*(19)+in_buf[325]*(21)+in_buf[326]*(8)+in_buf[327]*(5)+in_buf[328]*(24)+in_buf[329]*(17)+in_buf[330]*(22)+in_buf[331]*(23)+in_buf[332]*(34)+in_buf[333]*(32)+in_buf[334]*(33)+in_buf[335]*(25)+in_buf[336]*(6)+in_buf[337]*(0)+in_buf[338]*(39)+in_buf[339]*(44)+in_buf[340]*(23)+in_buf[341]*(5)+in_buf[342]*(8)+in_buf[343]*(-4)+in_buf[344]*(5)+in_buf[345]*(-1)+in_buf[346]*(-17)+in_buf[347]*(-9)+in_buf[348]*(-6)+in_buf[349]*(22)+in_buf[350]*(37)+in_buf[351]*(21)+in_buf[352]*(-2)+in_buf[353]*(6)+in_buf[354]*(2)+in_buf[355]*(9)+in_buf[356]*(12)+in_buf[357]*(15)+in_buf[358]*(7)+in_buf[359]*(10)+in_buf[360]*(-18)+in_buf[361]*(9)+in_buf[362]*(48)+in_buf[363]*(34)+in_buf[364]*(-17)+in_buf[365]*(-1)+in_buf[366]*(18)+in_buf[367]*(31)+in_buf[368]*(28)+in_buf[369]*(-13)+in_buf[370]*(-10)+in_buf[371]*(6)+in_buf[372]*(-5)+in_buf[373]*(-1)+in_buf[374]*(-9)+in_buf[375]*(-6)+in_buf[376]*(5)+in_buf[377]*(26)+in_buf[378]*(17)+in_buf[379]*(-3)+in_buf[380]*(-2)+in_buf[381]*(-4)+in_buf[382]*(-10)+in_buf[383]*(0)+in_buf[384]*(4)+in_buf[385]*(9)+in_buf[386]*(9)+in_buf[387]*(0)+in_buf[388]*(-25)+in_buf[389]*(1)+in_buf[390]*(30)+in_buf[391]*(1)+in_buf[392]*(0)+in_buf[393]*(-4)+in_buf[394]*(-4)+in_buf[395]*(19)+in_buf[396]*(8)+in_buf[397]*(-18)+in_buf[398]*(-10)+in_buf[399]*(-2)+in_buf[400]*(-1)+in_buf[401]*(-6)+in_buf[402]*(-6)+in_buf[403]*(-1)+in_buf[404]*(9)+in_buf[405]*(8)+in_buf[406]*(-11)+in_buf[407]*(-12)+in_buf[408]*(-2)+in_buf[409]*(-3)+in_buf[410]*(4)+in_buf[411]*(6)+in_buf[412]*(8)+in_buf[413]*(0)+in_buf[414]*(-4)+in_buf[415]*(-2)+in_buf[416]*(11)+in_buf[417]*(-7)+in_buf[418]*(0)+in_buf[419]*(6)+in_buf[420]*(-3)+in_buf[421]*(-1)+in_buf[422]*(-28)+in_buf[423]*(-9)+in_buf[424]*(8)+in_buf[425]*(16)+in_buf[426]*(10)+in_buf[427]*(0)+in_buf[428]*(7)+in_buf[429]*(4)+in_buf[430]*(3)+in_buf[431]*(15)+in_buf[432]*(3)+in_buf[433]*(-17)+in_buf[434]*(-30)+in_buf[435]*(-20)+in_buf[436]*(-3)+in_buf[437]*(7)+in_buf[438]*(14)+in_buf[439]*(7)+in_buf[440]*(12)+in_buf[441]*(-7)+in_buf[442]*(-10)+in_buf[443]*(9)+in_buf[444]*(15)+in_buf[445]*(1)+in_buf[446]*(4)+in_buf[447]*(-14)+in_buf[448]*(-14)+in_buf[449]*(-13)+in_buf[450]*(-10)+in_buf[451]*(-7)+in_buf[452]*(19)+in_buf[453]*(23)+in_buf[454]*(14)+in_buf[455]*(-2)+in_buf[456]*(10)+in_buf[457]*(-8)+in_buf[458]*(-1)+in_buf[459]*(12)+in_buf[460]*(6)+in_buf[461]*(-13)+in_buf[462]*(-29)+in_buf[463]*(-19)+in_buf[464]*(-3)+in_buf[465]*(3)+in_buf[466]*(10)+in_buf[467]*(2)+in_buf[468]*(-2)+in_buf[469]*(-25)+in_buf[470]*(-8)+in_buf[471]*(10)+in_buf[472]*(6)+in_buf[473]*(-4)+in_buf[474]*(-12)+in_buf[475]*(0)+in_buf[476]*(-2)+in_buf[477]*(9)+in_buf[478]*(-29)+in_buf[479]*(4)+in_buf[480]*(11)+in_buf[481]*(24)+in_buf[482]*(18)+in_buf[483]*(1)+in_buf[484]*(11)+in_buf[485]*(4)+in_buf[486]*(2)+in_buf[487]*(-5)+in_buf[488]*(-2)+in_buf[489]*(1)+in_buf[490]*(-1)+in_buf[491]*(6)+in_buf[492]*(0)+in_buf[493]*(8)+in_buf[494]*(4)+in_buf[495]*(12)+in_buf[496]*(11)+in_buf[497]*(-16)+in_buf[498]*(-6)+in_buf[499]*(0)+in_buf[500]*(19)+in_buf[501]*(8)+in_buf[502]*(-5)+in_buf[503]*(16)+in_buf[504]*(35)+in_buf[505]*(9)+in_buf[506]*(-19)+in_buf[507]*(-17)+in_buf[508]*(2)+in_buf[509]*(12)+in_buf[510]*(18)+in_buf[511]*(16)+in_buf[512]*(16)+in_buf[513]*(8)+in_buf[514]*(8)+in_buf[515]*(9)+in_buf[516]*(9)+in_buf[517]*(10)+in_buf[518]*(0)+in_buf[519]*(-3)+in_buf[520]*(-11)+in_buf[521]*(8)+in_buf[522]*(1)+in_buf[523]*(7)+in_buf[524]*(13)+in_buf[525]*(-10)+in_buf[526]*(2)+in_buf[527]*(-2)+in_buf[528]*(0)+in_buf[529]*(5)+in_buf[530]*(3)+in_buf[531]*(-22)+in_buf[532]*(-6)+in_buf[533]*(36)+in_buf[534]*(11)+in_buf[535]*(-24)+in_buf[536]*(-11)+in_buf[537]*(7)+in_buf[538]*(22)+in_buf[539]*(14)+in_buf[540]*(11)+in_buf[541]*(13)+in_buf[542]*(5)+in_buf[543]*(0)+in_buf[544]*(17)+in_buf[545]*(-1)+in_buf[546]*(-19)+in_buf[547]*(-17)+in_buf[548]*(-14)+in_buf[549]*(-3)+in_buf[550]*(4)+in_buf[551]*(1)+in_buf[552]*(0)+in_buf[553]*(-13)+in_buf[554]*(-10)+in_buf[555]*(-8)+in_buf[556]*(20)+in_buf[557]*(16)+in_buf[558]*(-29)+in_buf[559]*(-1)+in_buf[560]*(0)+in_buf[561]*(27)+in_buf[562]*(-24)+in_buf[563]*(-53)+in_buf[564]*(-12)+in_buf[565]*(12)+in_buf[566]*(7)+in_buf[567]*(-24)+in_buf[568]*(6)+in_buf[569]*(8)+in_buf[570]*(-5)+in_buf[571]*(-17)+in_buf[572]*(-12)+in_buf[573]*(-8)+in_buf[574]*(-33)+in_buf[575]*(-27)+in_buf[576]*(-10)+in_buf[577]*(10)+in_buf[578]*(-1)+in_buf[579]*(1)+in_buf[580]*(-15)+in_buf[581]*(-12)+in_buf[582]*(-7)+in_buf[583]*(-1)+in_buf[584]*(28)+in_buf[585]*(36)+in_buf[586]*(-37)+in_buf[587]*(7)+in_buf[588]*(-9)+in_buf[589]*(1)+in_buf[590]*(-35)+in_buf[591]*(-42)+in_buf[592]*(-16)+in_buf[593]*(-4)+in_buf[594]*(-12)+in_buf[595]*(-25)+in_buf[596]*(-28)+in_buf[597]*(-16)+in_buf[598]*(-14)+in_buf[599]*(-33)+in_buf[600]*(-16)+in_buf[601]*(-31)+in_buf[602]*(-34)+in_buf[603]*(-13)+in_buf[604]*(0)+in_buf[605]*(-2)+in_buf[606]*(1)+in_buf[607]*(-6)+in_buf[608]*(10)+in_buf[609]*(7)+in_buf[610]*(-21)+in_buf[611]*(-7)+in_buf[612]*(31)+in_buf[613]*(31)+in_buf[614]*(-2)+in_buf[615]*(3)+in_buf[616]*(-13)+in_buf[617]*(-7)+in_buf[618]*(-37)+in_buf[619]*(3)+in_buf[620]*(-3)+in_buf[621]*(-12)+in_buf[622]*(-15)+in_buf[623]*(-25)+in_buf[624]*(-15)+in_buf[625]*(-10)+in_buf[626]*(-21)+in_buf[627]*(-19)+in_buf[628]*(-6)+in_buf[629]*(-7)+in_buf[630]*(-1)+in_buf[631]*(-7)+in_buf[632]*(12)+in_buf[633]*(5)+in_buf[634]*(-9)+in_buf[635]*(-15)+in_buf[636]*(0)+in_buf[637]*(-19)+in_buf[638]*(-15)+in_buf[639]*(21)+in_buf[640]*(28)+in_buf[641]*(23)+in_buf[642]*(22)+in_buf[643]*(10)+in_buf[644]*(4)+in_buf[645]*(2)+in_buf[646]*(-48)+in_buf[647]*(20)+in_buf[648]*(3)+in_buf[649]*(-6)+in_buf[650]*(-21)+in_buf[651]*(-23)+in_buf[652]*(0)+in_buf[653]*(-3)+in_buf[654]*(-1)+in_buf[655]*(3)+in_buf[656]*(20)+in_buf[657]*(16)+in_buf[658]*(12)+in_buf[659]*(7)+in_buf[660]*(17)+in_buf[661]*(0)+in_buf[662]*(-21)+in_buf[663]*(-19)+in_buf[664]*(1)+in_buf[665]*(-17)+in_buf[666]*(2)+in_buf[667]*(37)+in_buf[668]*(32)+in_buf[669]*(16)+in_buf[670]*(4)+in_buf[671]*(-2)+in_buf[672]*(0)+in_buf[673]*(1)+in_buf[674]*(-13)+in_buf[675]*(10)+in_buf[676]*(19)+in_buf[677]*(23)+in_buf[678]*(-5)+in_buf[679]*(-2)+in_buf[680]*(0)+in_buf[681]*(-14)+in_buf[682]*(14)+in_buf[683]*(3)+in_buf[684]*(11)+in_buf[685]*(13)+in_buf[686]*(-2)+in_buf[687]*(13)+in_buf[688]*(-1)+in_buf[689]*(-15)+in_buf[690]*(-24)+in_buf[691]*(-8)+in_buf[692]*(3)+in_buf[693]*(-18)+in_buf[694]*(1)+in_buf[695]*(43)+in_buf[696]*(5)+in_buf[697]*(-17)+in_buf[698]*(-11)+in_buf[699]*(1)+in_buf[700]*(3)+in_buf[701]*(3)+in_buf[702]*(22)+in_buf[703]*(16)+in_buf[704]*(15)+in_buf[705]*(27)+in_buf[706]*(-5)+in_buf[707]*(3)+in_buf[708]*(0)+in_buf[709]*(9)+in_buf[710]*(2)+in_buf[711]*(10)+in_buf[712]*(4)+in_buf[713]*(13)+in_buf[714]*(12)+in_buf[715]*(9)+in_buf[716]*(12)+in_buf[717]*(-5)+in_buf[718]*(-15)+in_buf[719]*(31)+in_buf[720]*(23)+in_buf[721]*(22)+in_buf[722]*(12)+in_buf[723]*(15)+in_buf[724]*(31)+in_buf[725]*(0)+in_buf[726]*(-11)+in_buf[727]*(4)+in_buf[728]*(2)+in_buf[729]*(4)+in_buf[730]*(-2)+in_buf[731]*(23)+in_buf[732]*(14)+in_buf[733]*(29)+in_buf[734]*(32)+in_buf[735]*(28)+in_buf[736]*(26)+in_buf[737]*(47)+in_buf[738]*(24)+in_buf[739]*(24)+in_buf[740]*(41)+in_buf[741]*(57)+in_buf[742]*(71)+in_buf[743]*(22)+in_buf[744]*(33)+in_buf[745]*(35)+in_buf[746]*(33)+in_buf[747]*(48)+in_buf[748]*(72)+in_buf[749]*(52)+in_buf[750]*(52)+in_buf[751]*(4)+in_buf[752]*(13)+in_buf[753]*(-1)+in_buf[754]*(-3)+in_buf[755]*(2)+in_buf[756]*(0)+in_buf[757]*(2)+in_buf[758]*(-2)+in_buf[759]*(1)+in_buf[760]*(-24)+in_buf[761]*(-14)+in_buf[762]*(13)+in_buf[763]*(18)+in_buf[764]*(17)+in_buf[765]*(9)+in_buf[766]*(47)+in_buf[767]*(37)+in_buf[768]*(28)+in_buf[769]*(-7)+in_buf[770]*(51)+in_buf[771]*(32)+in_buf[772]*(24)+in_buf[773]*(-3)+in_buf[774]*(4)+in_buf[775]*(38)+in_buf[776]*(16)+in_buf[777]*(22)+in_buf[778]*(19)+in_buf[779]*(-26)+in_buf[780]*(-1)+in_buf[781]*(0)+in_buf[782]*(0)+in_buf[783]*(0);
assign in_buf_weight035=in_buf[0]*(-3)+in_buf[1]*(1)+in_buf[2]*(-2)+in_buf[3]*(4)+in_buf[4]*(4)+in_buf[5]*(4)+in_buf[6]*(0)+in_buf[7]*(1)+in_buf[8]*(0)+in_buf[9]*(0)+in_buf[10]*(-2)+in_buf[11]*(-3)+in_buf[12]*(20)+in_buf[13]*(20)+in_buf[14]*(7)+in_buf[15]*(6)+in_buf[16]*(0)+in_buf[17]*(1)+in_buf[18]*(0)+in_buf[19]*(3)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(-2)+in_buf[23]*(3)+in_buf[24]*(-2)+in_buf[25]*(-3)+in_buf[26]*(0)+in_buf[27]*(-3)+in_buf[28]*(4)+in_buf[29]*(2)+in_buf[30]*(-2)+in_buf[31]*(-2)+in_buf[32]*(2)+in_buf[33]*(3)+in_buf[34]*(12)+in_buf[35]*(16)+in_buf[36]*(18)+in_buf[37]*(24)+in_buf[38]*(37)+in_buf[39]*(35)+in_buf[40]*(45)+in_buf[41]*(14)+in_buf[42]*(-9)+in_buf[43]*(52)+in_buf[44]*(39)+in_buf[45]*(62)+in_buf[46]*(39)+in_buf[47]*(32)+in_buf[48]*(32)+in_buf[49]*(25)+in_buf[50]*(21)+in_buf[51]*(10)+in_buf[52]*(0)+in_buf[53]*(0)+in_buf[54]*(-3)+in_buf[55]*(-2)+in_buf[56]*(1)+in_buf[57]*(-3)+in_buf[58]*(19)+in_buf[59]*(10)+in_buf[60]*(16)+in_buf[61]*(7)+in_buf[62]*(18)+in_buf[63]*(20)+in_buf[64]*(8)+in_buf[65]*(2)+in_buf[66]*(10)+in_buf[67]*(53)+in_buf[68]*(37)+in_buf[69]*(27)+in_buf[70]*(27)+in_buf[71]*(35)+in_buf[72]*(23)+in_buf[73]*(40)+in_buf[74]*(61)+in_buf[75]*(43)+in_buf[76]*(43)+in_buf[77]*(39)+in_buf[78]*(52)+in_buf[79]*(37)+in_buf[80]*(2)+in_buf[81]*(-5)+in_buf[82]*(4)+in_buf[83]*(2)+in_buf[84]*(2)+in_buf[85]*(2)+in_buf[86]*(15)+in_buf[87]*(8)+in_buf[88]*(-7)+in_buf[89]*(-14)+in_buf[90]*(11)+in_buf[91]*(-6)+in_buf[92]*(1)+in_buf[93]*(17)+in_buf[94]*(-7)+in_buf[95]*(16)+in_buf[96]*(20)+in_buf[97]*(32)+in_buf[98]*(22)+in_buf[99]*(15)+in_buf[100]*(16)+in_buf[101]*(-6)+in_buf[102]*(2)+in_buf[103]*(18)+in_buf[104]*(-2)+in_buf[105]*(7)+in_buf[106]*(1)+in_buf[107]*(12)+in_buf[108]*(-15)+in_buf[109]*(-17)+in_buf[110]*(0)+in_buf[111]*(4)+in_buf[112]*(0)+in_buf[113]*(1)+in_buf[114]*(21)+in_buf[115]*(-15)+in_buf[116]*(2)+in_buf[117]*(-38)+in_buf[118]*(-35)+in_buf[119]*(-42)+in_buf[120]*(-24)+in_buf[121]*(-16)+in_buf[122]*(-9)+in_buf[123]*(-8)+in_buf[124]*(-8)+in_buf[125]*(5)+in_buf[126]*(14)+in_buf[127]*(10)+in_buf[128]*(13)+in_buf[129]*(17)+in_buf[130]*(11)+in_buf[131]*(12)+in_buf[132]*(-14)+in_buf[133]*(-37)+in_buf[134]*(-44)+in_buf[135]*(-24)+in_buf[136]*(-46)+in_buf[137]*(-39)+in_buf[138]*(-11)+in_buf[139]*(1)+in_buf[140]*(0)+in_buf[141]*(-1)+in_buf[142]*(54)+in_buf[143]*(-27)+in_buf[144]*(-35)+in_buf[145]*(-34)+in_buf[146]*(-35)+in_buf[147]*(-27)+in_buf[148]*(-10)+in_buf[149]*(-30)+in_buf[150]*(-16)+in_buf[151]*(-4)+in_buf[152]*(0)+in_buf[153]*(3)+in_buf[154]*(13)+in_buf[155]*(14)+in_buf[156]*(2)+in_buf[157]*(-4)+in_buf[158]*(-4)+in_buf[159]*(-12)+in_buf[160]*(-29)+in_buf[161]*(-31)+in_buf[162]*(-39)+in_buf[163]*(-25)+in_buf[164]*(-38)+in_buf[165]*(-28)+in_buf[166]*(-9)+in_buf[167]*(3)+in_buf[168]*(0)+in_buf[169]*(-16)+in_buf[170]*(-14)+in_buf[171]*(-20)+in_buf[172]*(-29)+in_buf[173]*(-36)+in_buf[174]*(-34)+in_buf[175]*(-33)+in_buf[176]*(-34)+in_buf[177]*(-30)+in_buf[178]*(-8)+in_buf[179]*(17)+in_buf[180]*(17)+in_buf[181]*(22)+in_buf[182]*(37)+in_buf[183]*(26)+in_buf[184]*(28)+in_buf[185]*(14)+in_buf[186]*(-13)+in_buf[187]*(-39)+in_buf[188]*(-45)+in_buf[189]*(-30)+in_buf[190]*(-34)+in_buf[191]*(-46)+in_buf[192]*(-39)+in_buf[193]*(-7)+in_buf[194]*(11)+in_buf[195]*(0)+in_buf[196]*(0)+in_buf[197]*(-14)+in_buf[198]*(-5)+in_buf[199]*(-10)+in_buf[200]*(-36)+in_buf[201]*(-44)+in_buf[202]*(-32)+in_buf[203]*(-39)+in_buf[204]*(-26)+in_buf[205]*(-17)+in_buf[206]*(3)+in_buf[207]*(17)+in_buf[208]*(31)+in_buf[209]*(27)+in_buf[210]*(35)+in_buf[211]*(43)+in_buf[212]*(26)+in_buf[213]*(-8)+in_buf[214]*(-17)+in_buf[215]*(-39)+in_buf[216]*(-36)+in_buf[217]*(-18)+in_buf[218]*(-27)+in_buf[219]*(-45)+in_buf[220]*(-28)+in_buf[221]*(-14)+in_buf[222]*(1)+in_buf[223]*(-23)+in_buf[224]*(4)+in_buf[225]*(-6)+in_buf[226]*(0)+in_buf[227]*(2)+in_buf[228]*(-14)+in_buf[229]*(-18)+in_buf[230]*(-9)+in_buf[231]*(-29)+in_buf[232]*(8)+in_buf[233]*(-1)+in_buf[234]*(3)+in_buf[235]*(15)+in_buf[236]*(8)+in_buf[237]*(17)+in_buf[238]*(26)+in_buf[239]*(15)+in_buf[240]*(-14)+in_buf[241]*(-33)+in_buf[242]*(-31)+in_buf[243]*(-14)+in_buf[244]*(-21)+in_buf[245]*(-10)+in_buf[246]*(-37)+in_buf[247]*(-51)+in_buf[248]*(-38)+in_buf[249]*(-18)+in_buf[250]*(5)+in_buf[251]*(-14)+in_buf[252]*(1)+in_buf[253]*(-11)+in_buf[254]*(8)+in_buf[255]*(29)+in_buf[256]*(-1)+in_buf[257]*(0)+in_buf[258]*(-2)+in_buf[259]*(4)+in_buf[260]*(4)+in_buf[261]*(12)+in_buf[262]*(12)+in_buf[263]*(3)+in_buf[264]*(6)+in_buf[265]*(28)+in_buf[266]*(31)+in_buf[267]*(-5)+in_buf[268]*(-28)+in_buf[269]*(-35)+in_buf[270]*(-33)+in_buf[271]*(-19)+in_buf[272]*(-3)+in_buf[273]*(-8)+in_buf[274]*(-41)+in_buf[275]*(-41)+in_buf[276]*(-7)+in_buf[277]*(-12)+in_buf[278]*(-9)+in_buf[279]*(-3)+in_buf[280]*(2)+in_buf[281]*(-4)+in_buf[282]*(4)+in_buf[283]*(22)+in_buf[284]*(-17)+in_buf[285]*(6)+in_buf[286]*(18)+in_buf[287]*(5)+in_buf[288]*(3)+in_buf[289]*(8)+in_buf[290]*(7)+in_buf[291]*(7)+in_buf[292]*(16)+in_buf[293]*(21)+in_buf[294]*(17)+in_buf[295]*(-15)+in_buf[296]*(-33)+in_buf[297]*(-29)+in_buf[298]*(-24)+in_buf[299]*(-11)+in_buf[300]*(-6)+in_buf[301]*(5)+in_buf[302]*(-14)+in_buf[303]*(7)+in_buf[304]*(-5)+in_buf[305]*(-27)+in_buf[306]*(-15)+in_buf[307]*(-17)+in_buf[308]*(0)+in_buf[309]*(-16)+in_buf[310]*(-4)+in_buf[311]*(3)+in_buf[312]*(-7)+in_buf[313]*(2)+in_buf[314]*(23)+in_buf[315]*(13)+in_buf[316]*(5)+in_buf[317]*(18)+in_buf[318]*(5)+in_buf[319]*(-1)+in_buf[320]*(8)+in_buf[321]*(0)+in_buf[322]*(-6)+in_buf[323]*(-31)+in_buf[324]*(-19)+in_buf[325]*(-5)+in_buf[326]*(-8)+in_buf[327]*(3)+in_buf[328]*(6)+in_buf[329]*(28)+in_buf[330]*(29)+in_buf[331]*(20)+in_buf[332]*(10)+in_buf[333]*(3)+in_buf[334]*(1)+in_buf[335]*(-4)+in_buf[336]*(3)+in_buf[337]*(-2)+in_buf[338]*(22)+in_buf[339]*(-5)+in_buf[340]*(22)+in_buf[341]*(7)+in_buf[342]*(17)+in_buf[343]*(25)+in_buf[344]*(16)+in_buf[345]*(24)+in_buf[346]*(-5)+in_buf[347]*(-4)+in_buf[348]*(-24)+in_buf[349]*(-17)+in_buf[350]*(-9)+in_buf[351]*(-14)+in_buf[352]*(-3)+in_buf[353]*(6)+in_buf[354]*(-1)+in_buf[355]*(0)+in_buf[356]*(6)+in_buf[357]*(16)+in_buf[358]*(37)+in_buf[359]*(14)+in_buf[360]*(7)+in_buf[361]*(-23)+in_buf[362]*(-23)+in_buf[363]*(1)+in_buf[364]*(11)+in_buf[365]*(-1)+in_buf[366]*(-7)+in_buf[367]*(-5)+in_buf[368]*(9)+in_buf[369]*(-1)+in_buf[370]*(21)+in_buf[371]*(28)+in_buf[372]*(27)+in_buf[373]*(18)+in_buf[374]*(15)+in_buf[375]*(-2)+in_buf[376]*(-23)+in_buf[377]*(-25)+in_buf[378]*(-4)+in_buf[379]*(1)+in_buf[380]*(5)+in_buf[381]*(-6)+in_buf[382]*(-5)+in_buf[383]*(-3)+in_buf[384]*(-18)+in_buf[385]*(8)+in_buf[386]*(20)+in_buf[387]*(23)+in_buf[388]*(9)+in_buf[389]*(16)+in_buf[390]*(-5)+in_buf[391]*(14)+in_buf[392]*(-23)+in_buf[393]*(-15)+in_buf[394]*(-11)+in_buf[395]*(-2)+in_buf[396]*(-4)+in_buf[397]*(-20)+in_buf[398]*(3)+in_buf[399]*(20)+in_buf[400]*(14)+in_buf[401]*(5)+in_buf[402]*(12)+in_buf[403]*(1)+in_buf[404]*(-26)+in_buf[405]*(-13)+in_buf[406]*(-3)+in_buf[407]*(8)+in_buf[408]*(9)+in_buf[409]*(-2)+in_buf[410]*(14)+in_buf[411]*(0)+in_buf[412]*(1)+in_buf[413]*(18)+in_buf[414]*(31)+in_buf[415]*(6)+in_buf[416]*(-6)+in_buf[417]*(33)+in_buf[418]*(-10)+in_buf[419]*(7)+in_buf[420]*(-14)+in_buf[421]*(-10)+in_buf[422]*(-10)+in_buf[423]*(-14)+in_buf[424]*(-21)+in_buf[425]*(-22)+in_buf[426]*(-11)+in_buf[427]*(8)+in_buf[428]*(7)+in_buf[429]*(3)+in_buf[430]*(11)+in_buf[431]*(3)+in_buf[432]*(3)+in_buf[433]*(3)+in_buf[434]*(8)+in_buf[435]*(0)+in_buf[436]*(5)+in_buf[437]*(2)+in_buf[438]*(7)+in_buf[439]*(-2)+in_buf[440]*(-1)+in_buf[441]*(6)+in_buf[442]*(-6)+in_buf[443]*(-23)+in_buf[444]*(-12)+in_buf[445]*(30)+in_buf[446]*(-34)+in_buf[447]*(-2)+in_buf[448]*(6)+in_buf[449]*(-9)+in_buf[450]*(-11)+in_buf[451]*(-4)+in_buf[452]*(-3)+in_buf[453]*(-3)+in_buf[454]*(-6)+in_buf[455]*(-3)+in_buf[456]*(3)+in_buf[457]*(-5)+in_buf[458]*(12)+in_buf[459]*(21)+in_buf[460]*(3)+in_buf[461]*(-9)+in_buf[462]*(17)+in_buf[463]*(0)+in_buf[464]*(8)+in_buf[465]*(-3)+in_buf[466]*(-2)+in_buf[467]*(-20)+in_buf[468]*(-10)+in_buf[469]*(-2)+in_buf[470]*(0)+in_buf[471]*(-5)+in_buf[472]*(-2)+in_buf[473]*(47)+in_buf[474]*(-11)+in_buf[475]*(-14)+in_buf[476]*(4)+in_buf[477]*(-6)+in_buf[478]*(-8)+in_buf[479]*(-2)+in_buf[480]*(0)+in_buf[481]*(-8)+in_buf[482]*(-21)+in_buf[483]*(-4)+in_buf[484]*(1)+in_buf[485]*(-11)+in_buf[486]*(6)+in_buf[487]*(0)+in_buf[488]*(-4)+in_buf[489]*(0)+in_buf[490]*(20)+in_buf[491]*(9)+in_buf[492]*(3)+in_buf[493]*(-13)+in_buf[494]*(-14)+in_buf[495]*(-29)+in_buf[496]*(-4)+in_buf[497]*(-5)+in_buf[498]*(11)+in_buf[499]*(2)+in_buf[500]*(20)+in_buf[501]*(63)+in_buf[502]*(-4)+in_buf[503]*(27)+in_buf[504]*(-11)+in_buf[505]*(-1)+in_buf[506]*(-12)+in_buf[507]*(-8)+in_buf[508]*(-13)+in_buf[509]*(-29)+in_buf[510]*(-21)+in_buf[511]*(6)+in_buf[512]*(2)+in_buf[513]*(-8)+in_buf[514]*(-2)+in_buf[515]*(-21)+in_buf[516]*(-16)+in_buf[517]*(-3)+in_buf[518]*(13)+in_buf[519]*(13)+in_buf[520]*(-11)+in_buf[521]*(-9)+in_buf[522]*(-1)+in_buf[523]*(-16)+in_buf[524]*(-5)+in_buf[525]*(-3)+in_buf[526]*(12)+in_buf[527]*(9)+in_buf[528]*(19)+in_buf[529]*(65)+in_buf[530]*(-15)+in_buf[531]*(-13)+in_buf[532]*(5)+in_buf[533]*(-18)+in_buf[534]*(-7)+in_buf[535]*(-28)+in_buf[536]*(-28)+in_buf[537]*(-26)+in_buf[538]*(-23)+in_buf[539]*(10)+in_buf[540]*(7)+in_buf[541]*(5)+in_buf[542]*(-7)+in_buf[543]*(-17)+in_buf[544]*(-7)+in_buf[545]*(5)+in_buf[546]*(13)+in_buf[547]*(20)+in_buf[548]*(4)+in_buf[549]*(-2)+in_buf[550]*(-2)+in_buf[551]*(-7)+in_buf[552]*(-7)+in_buf[553]*(4)+in_buf[554]*(12)+in_buf[555]*(28)+in_buf[556]*(31)+in_buf[557]*(50)+in_buf[558]*(2)+in_buf[559]*(-12)+in_buf[560]*(4)+in_buf[561]*(7)+in_buf[562]*(7)+in_buf[563]*(-35)+in_buf[564]*(-24)+in_buf[565]*(-28)+in_buf[566]*(-9)+in_buf[567]*(-3)+in_buf[568]*(-11)+in_buf[569]*(1)+in_buf[570]*(11)+in_buf[571]*(17)+in_buf[572]*(30)+in_buf[573]*(19)+in_buf[574]*(31)+in_buf[575]*(17)+in_buf[576]*(0)+in_buf[577]*(-6)+in_buf[578]*(16)+in_buf[579]*(-1)+in_buf[580]*(0)+in_buf[581]*(16)+in_buf[582]*(20)+in_buf[583]*(22)+in_buf[584]*(31)+in_buf[585]*(30)+in_buf[586]*(7)+in_buf[587]*(-1)+in_buf[588]*(9)+in_buf[589]*(0)+in_buf[590]*(2)+in_buf[591]*(0)+in_buf[592]*(-3)+in_buf[593]*(-9)+in_buf[594]*(17)+in_buf[595]*(7)+in_buf[596]*(-3)+in_buf[597]*(15)+in_buf[598]*(27)+in_buf[599]*(30)+in_buf[600]*(37)+in_buf[601]*(25)+in_buf[602]*(24)+in_buf[603]*(6)+in_buf[604]*(-3)+in_buf[605]*(10)+in_buf[606]*(15)+in_buf[607]*(-5)+in_buf[608]*(-14)+in_buf[609]*(-19)+in_buf[610]*(-10)+in_buf[611]*(6)+in_buf[612]*(3)+in_buf[613]*(1)+in_buf[614]*(22)+in_buf[615]*(-1)+in_buf[616]*(8)+in_buf[617]*(8)+in_buf[618]*(-12)+in_buf[619]*(6)+in_buf[620]*(20)+in_buf[621]*(15)+in_buf[622]*(14)+in_buf[623]*(8)+in_buf[624]*(13)+in_buf[625]*(27)+in_buf[626]*(22)+in_buf[627]*(10)+in_buf[628]*(15)+in_buf[629]*(10)+in_buf[630]*(-8)+in_buf[631]*(-6)+in_buf[632]*(-7)+in_buf[633]*(-7)+in_buf[634]*(-2)+in_buf[635]*(-29)+in_buf[636]*(-22)+in_buf[637]*(-42)+in_buf[638]*(-17)+in_buf[639]*(-16)+in_buf[640]*(-15)+in_buf[641]*(9)+in_buf[642]*(-19)+in_buf[643]*(3)+in_buf[644]*(2)+in_buf[645]*(-2)+in_buf[646]*(-19)+in_buf[647]*(-14)+in_buf[648]*(-5)+in_buf[649]*(24)+in_buf[650]*(6)+in_buf[651]*(-18)+in_buf[652]*(-13)+in_buf[653]*(3)+in_buf[654]*(-5)+in_buf[655]*(-14)+in_buf[656]*(2)+in_buf[657]*(-10)+in_buf[658]*(-6)+in_buf[659]*(-1)+in_buf[660]*(3)+in_buf[661]*(1)+in_buf[662]*(-12)+in_buf[663]*(-9)+in_buf[664]*(-6)+in_buf[665]*(-17)+in_buf[666]*(-8)+in_buf[667]*(-2)+in_buf[668]*(-17)+in_buf[669]*(-11)+in_buf[670]*(-20)+in_buf[671]*(2)+in_buf[672]*(1)+in_buf[673]*(3)+in_buf[674]*(-16)+in_buf[675]*(-26)+in_buf[676]*(-19)+in_buf[677]*(6)+in_buf[678]*(-20)+in_buf[679]*(-27)+in_buf[680]*(-26)+in_buf[681]*(-14)+in_buf[682]*(0)+in_buf[683]*(-31)+in_buf[684]*(-33)+in_buf[685]*(-27)+in_buf[686]*(-17)+in_buf[687]*(4)+in_buf[688]*(1)+in_buf[689]*(6)+in_buf[690]*(17)+in_buf[691]*(10)+in_buf[692]*(-2)+in_buf[693]*(-6)+in_buf[694]*(-6)+in_buf[695]*(14)+in_buf[696]*(9)+in_buf[697]*(41)+in_buf[698]*(26)+in_buf[699]*(3)+in_buf[700]*(-1)+in_buf[701]*(-3)+in_buf[702]*(18)+in_buf[703]*(-2)+in_buf[704]*(-3)+in_buf[705]*(-16)+in_buf[706]*(-28)+in_buf[707]*(-42)+in_buf[708]*(-21)+in_buf[709]*(-15)+in_buf[710]*(-10)+in_buf[711]*(-25)+in_buf[712]*(-13)+in_buf[713]*(-6)+in_buf[714]*(11)+in_buf[715]*(-13)+in_buf[716]*(-7)+in_buf[717]*(15)+in_buf[718]*(25)+in_buf[719]*(22)+in_buf[720]*(18)+in_buf[721]*(20)+in_buf[722]*(-8)+in_buf[723]*(-16)+in_buf[724]*(-14)+in_buf[725]*(26)+in_buf[726]*(21)+in_buf[727]*(-2)+in_buf[728]*(0)+in_buf[729]*(3)+in_buf[730]*(-2)+in_buf[731]*(15)+in_buf[732]*(23)+in_buf[733]*(5)+in_buf[734]*(14)+in_buf[735]*(35)+in_buf[736]*(47)+in_buf[737]*(26)+in_buf[738]*(27)+in_buf[739]*(19)+in_buf[740]*(15)+in_buf[741]*(16)+in_buf[742]*(50)+in_buf[743]*(33)+in_buf[744]*(48)+in_buf[745]*(47)+in_buf[746]*(51)+in_buf[747]*(33)+in_buf[748]*(27)+in_buf[749]*(17)+in_buf[750]*(24)+in_buf[751]*(44)+in_buf[752]*(5)+in_buf[753]*(4)+in_buf[754]*(1)+in_buf[755]*(-3)+in_buf[756]*(4)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(-2)+in_buf[760]*(0)+in_buf[761]*(-10)+in_buf[762]*(0)+in_buf[763]*(9)+in_buf[764]*(4)+in_buf[765]*(21)+in_buf[766]*(46)+in_buf[767]*(37)+in_buf[768]*(41)+in_buf[769]*(52)+in_buf[770]*(78)+in_buf[771]*(63)+in_buf[772]*(51)+in_buf[773]*(43)+in_buf[774]*(44)+in_buf[775]*(62)+in_buf[776]*(36)+in_buf[777]*(6)+in_buf[778]*(5)+in_buf[779]*(8)+in_buf[780]*(1)+in_buf[781]*(3)+in_buf[782]*(-1)+in_buf[783]*(5);
assign in_buf_weight036=in_buf[0]*(4)+in_buf[1]*(0)+in_buf[2]*(4)+in_buf[3]*(0)+in_buf[4]*(2)+in_buf[5]*(1)+in_buf[6]*(2)+in_buf[7]*(-1)+in_buf[8]*(0)+in_buf[9]*(3)+in_buf[10]*(5)+in_buf[11]*(2)+in_buf[12]*(-6)+in_buf[13]*(-5)+in_buf[14]*(-3)+in_buf[15]*(0)+in_buf[16]*(0)+in_buf[17]*(3)+in_buf[18]*(1)+in_buf[19]*(4)+in_buf[20]*(-2)+in_buf[21]*(4)+in_buf[22]*(3)+in_buf[23]*(0)+in_buf[24]*(-3)+in_buf[25]*(-2)+in_buf[26]*(0)+in_buf[27]*(-1)+in_buf[28]*(-1)+in_buf[29]*(4)+in_buf[30]*(-2)+in_buf[31]*(4)+in_buf[32]*(0)+in_buf[33]*(-2)+in_buf[34]*(-5)+in_buf[35]*(-8)+in_buf[36]*(-6)+in_buf[37]*(-5)+in_buf[38]*(-5)+in_buf[39]*(-4)+in_buf[40]*(-15)+in_buf[41]*(-12)+in_buf[42]*(-8)+in_buf[43]*(-12)+in_buf[44]*(-5)+in_buf[45]*(-3)+in_buf[46]*(-9)+in_buf[47]*(-9)+in_buf[48]*(-10)+in_buf[49]*(-2)+in_buf[50]*(-8)+in_buf[51]*(-4)+in_buf[52]*(2)+in_buf[53]*(3)+in_buf[54]*(2)+in_buf[55]*(1)+in_buf[56]*(1)+in_buf[57]*(1)+in_buf[58]*(-5)+in_buf[59]*(2)+in_buf[60]*(1)+in_buf[61]*(-5)+in_buf[62]*(-7)+in_buf[63]*(-13)+in_buf[64]*(-11)+in_buf[65]*(-20)+in_buf[66]*(-9)+in_buf[67]*(-5)+in_buf[68]*(-29)+in_buf[69]*(-73)+in_buf[70]*(-74)+in_buf[71]*(-45)+in_buf[72]*(-33)+in_buf[73]*(3)+in_buf[74]*(8)+in_buf[75]*(6)+in_buf[76]*(9)+in_buf[77]*(-4)+in_buf[78]*(-6)+in_buf[79]*(-10)+in_buf[80]*(-1)+in_buf[81]*(0)+in_buf[82]*(1)+in_buf[83]*(0)+in_buf[84]*(3)+in_buf[85]*(-3)+in_buf[86]*(3)+in_buf[87]*(5)+in_buf[88]*(7)+in_buf[89]*(9)+in_buf[90]*(8)+in_buf[91]*(-14)+in_buf[92]*(-45)+in_buf[93]*(-49)+in_buf[94]*(-41)+in_buf[95]*(-5)+in_buf[96]*(-5)+in_buf[97]*(-23)+in_buf[98]*(-21)+in_buf[99]*(-9)+in_buf[100]*(-25)+in_buf[101]*(5)+in_buf[102]*(24)+in_buf[103]*(9)+in_buf[104]*(14)+in_buf[105]*(4)+in_buf[106]*(-10)+in_buf[107]*(-10)+in_buf[108]*(-29)+in_buf[109]*(-25)+in_buf[110]*(-26)+in_buf[111]*(0)+in_buf[112]*(-2)+in_buf[113]*(8)+in_buf[114]*(25)+in_buf[115]*(37)+in_buf[116]*(32)+in_buf[117]*(12)+in_buf[118]*(2)+in_buf[119]*(-3)+in_buf[120]*(-35)+in_buf[121]*(-34)+in_buf[122]*(-4)+in_buf[123]*(5)+in_buf[124]*(1)+in_buf[125]*(23)+in_buf[126]*(9)+in_buf[127]*(-3)+in_buf[128]*(-3)+in_buf[129]*(-4)+in_buf[130]*(13)+in_buf[131]*(10)+in_buf[132]*(4)+in_buf[133]*(5)+in_buf[134]*(15)+in_buf[135]*(20)+in_buf[136]*(13)+in_buf[137]*(-6)+in_buf[138]*(-16)+in_buf[139]*(-26)+in_buf[140]*(1)+in_buf[141]*(4)+in_buf[142]*(22)+in_buf[143]*(20)+in_buf[144]*(29)+in_buf[145]*(18)+in_buf[146]*(20)+in_buf[147]*(-6)+in_buf[148]*(-16)+in_buf[149]*(-6)+in_buf[150]*(5)+in_buf[151]*(6)+in_buf[152]*(6)+in_buf[153]*(6)+in_buf[154]*(-3)+in_buf[155]*(-12)+in_buf[156]*(3)+in_buf[157]*(8)+in_buf[158]*(-17)+in_buf[159]*(-8)+in_buf[160]*(-1)+in_buf[161]*(-3)+in_buf[162]*(13)+in_buf[163]*(6)+in_buf[164]*(0)+in_buf[165]*(10)+in_buf[166]*(-42)+in_buf[167]*(-12)+in_buf[168]*(3)+in_buf[169]*(23)+in_buf[170]*(13)+in_buf[171]*(3)+in_buf[172]*(-6)+in_buf[173]*(10)+in_buf[174]*(-3)+in_buf[175]*(-11)+in_buf[176]*(6)+in_buf[177]*(9)+in_buf[178]*(16)+in_buf[179]*(11)+in_buf[180]*(7)+in_buf[181]*(13)+in_buf[182]*(2)+in_buf[183]*(-20)+in_buf[184]*(-11)+in_buf[185]*(-7)+in_buf[186]*(-10)+in_buf[187]*(0)+in_buf[188]*(10)+in_buf[189]*(12)+in_buf[190]*(16)+in_buf[191]*(6)+in_buf[192]*(-5)+in_buf[193]*(-35)+in_buf[194]*(-29)+in_buf[195]*(-31)+in_buf[196]*(4)+in_buf[197]*(26)+in_buf[198]*(9)+in_buf[199]*(-20)+in_buf[200]*(-12)+in_buf[201]*(-13)+in_buf[202]*(-8)+in_buf[203]*(1)+in_buf[204]*(4)+in_buf[205]*(12)+in_buf[206]*(6)+in_buf[207]*(3)+in_buf[208]*(-4)+in_buf[209]*(-5)+in_buf[210]*(-2)+in_buf[211]*(-28)+in_buf[212]*(-17)+in_buf[213]*(0)+in_buf[214]*(6)+in_buf[215]*(15)+in_buf[216]*(14)+in_buf[217]*(-1)+in_buf[218]*(-3)+in_buf[219]*(12)+in_buf[220]*(11)+in_buf[221]*(-10)+in_buf[222]*(2)+in_buf[223]*(-24)+in_buf[224]*(-3)+in_buf[225]*(-18)+in_buf[226]*(22)+in_buf[227]*(14)+in_buf[228]*(5)+in_buf[229]*(6)+in_buf[230]*(0)+in_buf[231]*(11)+in_buf[232]*(0)+in_buf[233]*(2)+in_buf[234]*(-6)+in_buf[235]*(-11)+in_buf[236]*(1)+in_buf[237]*(2)+in_buf[238]*(-3)+in_buf[239]*(-11)+in_buf[240]*(-1)+in_buf[241]*(12)+in_buf[242]*(29)+in_buf[243]*(10)+in_buf[244]*(12)+in_buf[245]*(7)+in_buf[246]*(10)+in_buf[247]*(-5)+in_buf[248]*(23)+in_buf[249]*(16)+in_buf[250]*(4)+in_buf[251]*(0)+in_buf[252]*(-5)+in_buf[253]*(-14)+in_buf[254]*(33)+in_buf[255]*(26)+in_buf[256]*(8)+in_buf[257]*(-17)+in_buf[258]*(10)+in_buf[259]*(13)+in_buf[260]*(8)+in_buf[261]*(6)+in_buf[262]*(-6)+in_buf[263]*(-9)+in_buf[264]*(-8)+in_buf[265]*(-4)+in_buf[266]*(-8)+in_buf[267]*(-5)+in_buf[268]*(16)+in_buf[269]*(30)+in_buf[270]*(27)+in_buf[271]*(23)+in_buf[272]*(30)+in_buf[273]*(14)+in_buf[274]*(21)+in_buf[275]*(22)+in_buf[276]*(13)+in_buf[277]*(-22)+in_buf[278]*(-28)+in_buf[279]*(-48)+in_buf[280]*(-6)+in_buf[281]*(-4)+in_buf[282]*(17)+in_buf[283]*(26)+in_buf[284]*(35)+in_buf[285]*(-16)+in_buf[286]*(-24)+in_buf[287]*(-11)+in_buf[288]*(4)+in_buf[289]*(-8)+in_buf[290]*(-6)+in_buf[291]*(-22)+in_buf[292]*(-5)+in_buf[293]*(-17)+in_buf[294]*(-33)+in_buf[295]*(-5)+in_buf[296]*(1)+in_buf[297]*(10)+in_buf[298]*(11)+in_buf[299]*(10)+in_buf[300]*(21)+in_buf[301]*(5)+in_buf[302]*(18)+in_buf[303]*(44)+in_buf[304]*(10)+in_buf[305]*(12)+in_buf[306]*(-18)+in_buf[307]*(-37)+in_buf[308]*(-2)+in_buf[309]*(-5)+in_buf[310]*(-12)+in_buf[311]*(11)+in_buf[312]*(14)+in_buf[313]*(-1)+in_buf[314]*(-9)+in_buf[315]*(-19)+in_buf[316]*(-10)+in_buf[317]*(-6)+in_buf[318]*(0)+in_buf[319]*(-25)+in_buf[320]*(-11)+in_buf[321]*(-14)+in_buf[322]*(-17)+in_buf[323]*(3)+in_buf[324]*(0)+in_buf[325]*(0)+in_buf[326]*(-6)+in_buf[327]*(-10)+in_buf[328]*(1)+in_buf[329]*(0)+in_buf[330]*(23)+in_buf[331]*(22)+in_buf[332]*(35)+in_buf[333]*(32)+in_buf[334]*(4)+in_buf[335]*(-25)+in_buf[336]*(-1)+in_buf[337]*(1)+in_buf[338]*(6)+in_buf[339]*(-36)+in_buf[340]*(-3)+in_buf[341]*(-11)+in_buf[342]*(-6)+in_buf[343]*(-2)+in_buf[344]*(-13)+in_buf[345]*(-14)+in_buf[346]*(7)+in_buf[347]*(-2)+in_buf[348]*(3)+in_buf[349]*(22)+in_buf[350]*(0)+in_buf[351]*(0)+in_buf[352]*(0)+in_buf[353]*(-1)+in_buf[354]*(-9)+in_buf[355]*(-22)+in_buf[356]*(4)+in_buf[357]*(5)+in_buf[358]*(17)+in_buf[359]*(34)+in_buf[360]*(37)+in_buf[361]*(3)+in_buf[362]*(-42)+in_buf[363]*(-19)+in_buf[364]*(-11)+in_buf[365]*(4)+in_buf[366]*(-11)+in_buf[367]*(-37)+in_buf[368]*(-5)+in_buf[369]*(0)+in_buf[370]*(-2)+in_buf[371]*(16)+in_buf[372]*(12)+in_buf[373]*(23)+in_buf[374]*(22)+in_buf[375]*(11)+in_buf[376]*(19)+in_buf[377]*(10)+in_buf[378]*(0)+in_buf[379]*(6)+in_buf[380]*(0)+in_buf[381]*(-6)+in_buf[382]*(-17)+in_buf[383]*(-8)+in_buf[384]*(11)+in_buf[385]*(12)+in_buf[386]*(3)+in_buf[387]*(-1)+in_buf[388]*(-12)+in_buf[389]*(-23)+in_buf[390]*(-53)+in_buf[391]*(3)+in_buf[392]*(-10)+in_buf[393]*(7)+in_buf[394]*(-1)+in_buf[395]*(-20)+in_buf[396]*(-5)+in_buf[397]*(9)+in_buf[398]*(-10)+in_buf[399]*(11)+in_buf[400]*(30)+in_buf[401]*(37)+in_buf[402]*(24)+in_buf[403]*(21)+in_buf[404]*(37)+in_buf[405]*(21)+in_buf[406]*(19)+in_buf[407]*(18)+in_buf[408]*(4)+in_buf[409]*(15)+in_buf[410]*(0)+in_buf[411]*(-6)+in_buf[412]*(0)+in_buf[413]*(-9)+in_buf[414]*(-18)+in_buf[415]*(-18)+in_buf[416]*(-35)+in_buf[417]*(-39)+in_buf[418]*(-42)+in_buf[419]*(-4)+in_buf[420]*(-7)+in_buf[421]*(9)+in_buf[422]*(24)+in_buf[423]*(22)+in_buf[424]*(-9)+in_buf[425]*(-11)+in_buf[426]*(-21)+in_buf[427]*(-12)+in_buf[428]*(14)+in_buf[429]*(25)+in_buf[430]*(43)+in_buf[431]*(43)+in_buf[432]*(47)+in_buf[433]*(36)+in_buf[434]*(31)+in_buf[435]*(30)+in_buf[436]*(8)+in_buf[437]*(26)+in_buf[438]*(3)+in_buf[439]*(-11)+in_buf[440]*(-13)+in_buf[441]*(-23)+in_buf[442]*(7)+in_buf[443]*(-7)+in_buf[444]*(-38)+in_buf[445]*(-42)+in_buf[446]*(-18)+in_buf[447]*(5)+in_buf[448]*(-6)+in_buf[449]*(8)+in_buf[450]*(20)+in_buf[451]*(16)+in_buf[452]*(-1)+in_buf[453]*(-32)+in_buf[454]*(-32)+in_buf[455]*(-20)+in_buf[456]*(-19)+in_buf[457]*(0)+in_buf[458]*(12)+in_buf[459]*(35)+in_buf[460]*(59)+in_buf[461]*(59)+in_buf[462]*(40)+in_buf[463]*(24)+in_buf[464]*(15)+in_buf[465]*(11)+in_buf[466]*(2)+in_buf[467]*(-10)+in_buf[468]*(-13)+in_buf[469]*(-17)+in_buf[470]*(-31)+in_buf[471]*(-25)+in_buf[472]*(-44)+in_buf[473]*(-46)+in_buf[474]*(-50)+in_buf[475]*(-22)+in_buf[476]*(-2)+in_buf[477]*(15)+in_buf[478]*(9)+in_buf[479]*(-10)+in_buf[480]*(-13)+in_buf[481]*(-52)+in_buf[482]*(-55)+in_buf[483]*(-37)+in_buf[484]*(-55)+in_buf[485]*(-35)+in_buf[486]*(-28)+in_buf[487]*(-3)+in_buf[488]*(16)+in_buf[489]*(30)+in_buf[490]*(12)+in_buf[491]*(12)+in_buf[492]*(6)+in_buf[493]*(-5)+in_buf[494]*(-7)+in_buf[495]*(-19)+in_buf[496]*(-9)+in_buf[497]*(-3)+in_buf[498]*(-23)+in_buf[499]*(-9)+in_buf[500]*(-11)+in_buf[501]*(5)+in_buf[502]*(-11)+in_buf[503]*(-29)+in_buf[504]*(-24)+in_buf[505]*(8)+in_buf[506]*(15)+in_buf[507]*(-29)+in_buf[508]*(-30)+in_buf[509]*(-54)+in_buf[510]*(-53)+in_buf[511]*(-74)+in_buf[512]*(-83)+in_buf[513]*(-65)+in_buf[514]*(-48)+in_buf[515]*(-18)+in_buf[516]*(-14)+in_buf[517]*(4)+in_buf[518]*(2)+in_buf[519]*(-3)+in_buf[520]*(12)+in_buf[521]*(-6)+in_buf[522]*(-3)+in_buf[523]*(-21)+in_buf[524]*(-11)+in_buf[525]*(0)+in_buf[526]*(-17)+in_buf[527]*(-8)+in_buf[528]*(-2)+in_buf[529]*(13)+in_buf[530]*(27)+in_buf[531]*(0)+in_buf[532]*(11)+in_buf[533]*(-29)+in_buf[534]*(2)+in_buf[535]*(-1)+in_buf[536]*(-13)+in_buf[537]*(-28)+in_buf[538]*(-32)+in_buf[539]*(-46)+in_buf[540]*(-60)+in_buf[541]*(-57)+in_buf[542]*(-50)+in_buf[543]*(-37)+in_buf[544]*(-36)+in_buf[545]*(-20)+in_buf[546]*(-6)+in_buf[547]*(-2)+in_buf[548]*(10)+in_buf[549]*(1)+in_buf[550]*(0)+in_buf[551]*(-15)+in_buf[552]*(-10)+in_buf[553]*(1)+in_buf[554]*(-26)+in_buf[555]*(-27)+in_buf[556]*(-45)+in_buf[557]*(-7)+in_buf[558]*(-2)+in_buf[559]*(16)+in_buf[560]*(-4)+in_buf[561]*(18)+in_buf[562]*(17)+in_buf[563]*(20)+in_buf[564]*(18)+in_buf[565]*(0)+in_buf[566]*(-7)+in_buf[567]*(-9)+in_buf[568]*(-26)+in_buf[569]*(-28)+in_buf[570]*(-32)+in_buf[571]*(-24)+in_buf[572]*(-36)+in_buf[573]*(-15)+in_buf[574]*(-9)+in_buf[575]*(0)+in_buf[576]*(4)+in_buf[577]*(17)+in_buf[578]*(16)+in_buf[579]*(7)+in_buf[580]*(0)+in_buf[581]*(5)+in_buf[582]*(-15)+in_buf[583]*(-34)+in_buf[584]*(-46)+in_buf[585]*(-34)+in_buf[586]*(11)+in_buf[587]*(1)+in_buf[588]*(20)+in_buf[589]*(15)+in_buf[590]*(27)+in_buf[591]*(31)+in_buf[592]*(40)+in_buf[593]*(15)+in_buf[594]*(21)+in_buf[595]*(23)+in_buf[596]*(15)+in_buf[597]*(0)+in_buf[598]*(1)+in_buf[599]*(11)+in_buf[600]*(-7)+in_buf[601]*(-14)+in_buf[602]*(-14)+in_buf[603]*(-1)+in_buf[604]*(1)+in_buf[605]*(3)+in_buf[606]*(7)+in_buf[607]*(-10)+in_buf[608]*(-17)+in_buf[609]*(-22)+in_buf[610]*(-41)+in_buf[611]*(-20)+in_buf[612]*(-19)+in_buf[613]*(-6)+in_buf[614]*(-5)+in_buf[615]*(0)+in_buf[616]*(19)+in_buf[617]*(36)+in_buf[618]*(31)+in_buf[619]*(18)+in_buf[620]*(31)+in_buf[621]*(33)+in_buf[622]*(28)+in_buf[623]*(31)+in_buf[624]*(17)+in_buf[625]*(17)+in_buf[626]*(23)+in_buf[627]*(27)+in_buf[628]*(10)+in_buf[629]*(1)+in_buf[630]*(0)+in_buf[631]*(8)+in_buf[632]*(-4)+in_buf[633]*(-7)+in_buf[634]*(-4)+in_buf[635]*(2)+in_buf[636]*(-18)+in_buf[637]*(-37)+in_buf[638]*(-57)+in_buf[639]*(-26)+in_buf[640]*(-14)+in_buf[641]*(-2)+in_buf[642]*(27)+in_buf[643]*(-2)+in_buf[644]*(2)+in_buf[645]*(-3)+in_buf[646]*(30)+in_buf[647]*(25)+in_buf[648]*(40)+in_buf[649]*(36)+in_buf[650]*(24)+in_buf[651]*(28)+in_buf[652]*(25)+in_buf[653]*(19)+in_buf[654]*(28)+in_buf[655]*(21)+in_buf[656]*(3)+in_buf[657]*(8)+in_buf[658]*(12)+in_buf[659]*(4)+in_buf[660]*(-7)+in_buf[661]*(-9)+in_buf[662]*(-21)+in_buf[663]*(-32)+in_buf[664]*(-45)+in_buf[665]*(-61)+in_buf[666]*(-50)+in_buf[667]*(-21)+in_buf[668]*(-17)+in_buf[669]*(7)+in_buf[670]*(45)+in_buf[671]*(2)+in_buf[672]*(-3)+in_buf[673]*(-3)+in_buf[674]*(16)+in_buf[675]*(36)+in_buf[676]*(20)+in_buf[677]*(30)+in_buf[678]*(38)+in_buf[679]*(26)+in_buf[680]*(19)+in_buf[681]*(24)+in_buf[682]*(36)+in_buf[683]*(27)+in_buf[684]*(7)+in_buf[685]*(9)+in_buf[686]*(3)+in_buf[687]*(-17)+in_buf[688]*(-18)+in_buf[689]*(-33)+in_buf[690]*(-38)+in_buf[691]*(-43)+in_buf[692]*(-50)+in_buf[693]*(-28)+in_buf[694]*(-23)+in_buf[695]*(2)+in_buf[696]*(-14)+in_buf[697]*(7)+in_buf[698]*(-4)+in_buf[699]*(5)+in_buf[700]*(-3)+in_buf[701]*(4)+in_buf[702]*(10)+in_buf[703]*(-15)+in_buf[704]*(5)+in_buf[705]*(36)+in_buf[706]*(19)+in_buf[707]*(17)+in_buf[708]*(9)+in_buf[709]*(-4)+in_buf[710]*(15)+in_buf[711]*(5)+in_buf[712]*(10)+in_buf[713]*(7)+in_buf[714]*(-30)+in_buf[715]*(-36)+in_buf[716]*(-28)+in_buf[717]*(-40)+in_buf[718]*(-37)+in_buf[719]*(-25)+in_buf[720]*(-26)+in_buf[721]*(-11)+in_buf[722]*(18)+in_buf[723]*(26)+in_buf[724]*(6)+in_buf[725]*(7)+in_buf[726]*(-3)+in_buf[727]*(-3)+in_buf[728]*(-2)+in_buf[729]*(-1)+in_buf[730]*(3)+in_buf[731]*(-7)+in_buf[732]*(12)+in_buf[733]*(31)+in_buf[734]*(29)+in_buf[735]*(0)+in_buf[736]*(-22)+in_buf[737]*(-36)+in_buf[738]*(3)+in_buf[739]*(0)+in_buf[740]*(-18)+in_buf[741]*(-35)+in_buf[742]*(-31)+in_buf[743]*(-14)+in_buf[744]*(9)+in_buf[745]*(9)+in_buf[746]*(-23)+in_buf[747]*(-30)+in_buf[748]*(-25)+in_buf[749]*(0)+in_buf[750]*(-14)+in_buf[751]*(-2)+in_buf[752]*(28)+in_buf[753]*(-16)+in_buf[754]*(-2)+in_buf[755]*(-1)+in_buf[756]*(-1)+in_buf[757]*(4)+in_buf[758]*(-2)+in_buf[759]*(2)+in_buf[760]*(-27)+in_buf[761]*(-37)+in_buf[762]*(-35)+in_buf[763]*(-22)+in_buf[764]*(-20)+in_buf[765]*(-12)+in_buf[766]*(-36)+in_buf[767]*(-23)+in_buf[768]*(-9)+in_buf[769]*(-26)+in_buf[770]*(-9)+in_buf[771]*(4)+in_buf[772]*(-11)+in_buf[773]*(-25)+in_buf[774]*(-5)+in_buf[775]*(20)+in_buf[776]*(8)+in_buf[777]*(-6)+in_buf[778]*(-6)+in_buf[779]*(0)+in_buf[780]*(1)+in_buf[781]*(2)+in_buf[782]*(0)+in_buf[783]*(-1);
assign in_buf_weight037=in_buf[0]*(-3)+in_buf[1]*(4)+in_buf[2]*(-2)+in_buf[3]*(-2)+in_buf[4]*(1)+in_buf[5]*(4)+in_buf[6]*(0)+in_buf[7]*(0)+in_buf[8]*(-2)+in_buf[9]*(0)+in_buf[10]*(-2)+in_buf[11]*(1)+in_buf[12]*(-8)+in_buf[13]*(-11)+in_buf[14]*(4)+in_buf[15]*(0)+in_buf[16]*(-1)+in_buf[17]*(-1)+in_buf[18]*(-3)+in_buf[19]*(0)+in_buf[20]*(3)+in_buf[21]*(-1)+in_buf[22]*(3)+in_buf[23]*(4)+in_buf[24]*(1)+in_buf[25]*(-2)+in_buf[26]*(2)+in_buf[27]*(-2)+in_buf[28]*(4)+in_buf[29]*(0)+in_buf[30]*(2)+in_buf[31]*(0)+in_buf[32]*(-4)+in_buf[33]*(-4)+in_buf[34]*(-11)+in_buf[35]*(-10)+in_buf[36]*(-19)+in_buf[37]*(-12)+in_buf[38]*(-13)+in_buf[39]*(10)+in_buf[40]*(4)+in_buf[41]*(-4)+in_buf[42]*(-33)+in_buf[43]*(20)+in_buf[44]*(19)+in_buf[45]*(7)+in_buf[46]*(-27)+in_buf[47]*(-11)+in_buf[48]*(-13)+in_buf[49]*(-17)+in_buf[50]*(-4)+in_buf[51]*(-4)+in_buf[52]*(-2)+in_buf[53]*(0)+in_buf[54]*(4)+in_buf[55]*(2)+in_buf[56]*(3)+in_buf[57]*(-1)+in_buf[58]*(-19)+in_buf[59]*(8)+in_buf[60]*(4)+in_buf[61]*(-7)+in_buf[62]*(-21)+in_buf[63]*(-22)+in_buf[64]*(-17)+in_buf[65]*(-37)+in_buf[66]*(-51)+in_buf[67]*(-47)+in_buf[68]*(-16)+in_buf[69]*(-26)+in_buf[70]*(-48)+in_buf[71]*(-27)+in_buf[72]*(0)+in_buf[73]*(4)+in_buf[74]*(-28)+in_buf[75]*(-34)+in_buf[76]*(-33)+in_buf[77]*(-16)+in_buf[78]*(-19)+in_buf[79]*(-10)+in_buf[80]*(4)+in_buf[81]*(6)+in_buf[82]*(1)+in_buf[83]*(-3)+in_buf[84]*(2)+in_buf[85]*(-3)+in_buf[86]*(-19)+in_buf[87]*(-1)+in_buf[88]*(8)+in_buf[89]*(-7)+in_buf[90]*(-34)+in_buf[91]*(-7)+in_buf[92]*(-20)+in_buf[93]*(-24)+in_buf[94]*(-36)+in_buf[95]*(-25)+in_buf[96]*(-32)+in_buf[97]*(-38)+in_buf[98]*(-44)+in_buf[99]*(-23)+in_buf[100]*(-16)+in_buf[101]*(-9)+in_buf[102]*(-12)+in_buf[103]*(-28)+in_buf[104]*(-36)+in_buf[105]*(-22)+in_buf[106]*(-22)+in_buf[107]*(-32)+in_buf[108]*(6)+in_buf[109]*(11)+in_buf[110]*(8)+in_buf[111]*(4)+in_buf[112]*(0)+in_buf[113]*(-3)+in_buf[114]*(-7)+in_buf[115]*(29)+in_buf[116]*(1)+in_buf[117]*(-10)+in_buf[118]*(-9)+in_buf[119]*(-17)+in_buf[120]*(-37)+in_buf[121]*(-33)+in_buf[122]*(-50)+in_buf[123]*(-51)+in_buf[124]*(-60)+in_buf[125]*(-63)+in_buf[126]*(-82)+in_buf[127]*(-53)+in_buf[128]*(-50)+in_buf[129]*(-10)+in_buf[130]*(4)+in_buf[131]*(-16)+in_buf[132]*(-30)+in_buf[133]*(10)+in_buf[134]*(26)+in_buf[135]*(32)+in_buf[136]*(28)+in_buf[137]*(14)+in_buf[138]*(23)+in_buf[139]*(-15)+in_buf[140]*(-2)+in_buf[141]*(2)+in_buf[142]*(-27)+in_buf[143]*(5)+in_buf[144]*(-10)+in_buf[145]*(-6)+in_buf[146]*(-20)+in_buf[147]*(-26)+in_buf[148]*(-13)+in_buf[149]*(-12)+in_buf[150]*(-28)+in_buf[151]*(-21)+in_buf[152]*(-23)+in_buf[153]*(-22)+in_buf[154]*(-42)+in_buf[155]*(-45)+in_buf[156]*(-50)+in_buf[157]*(-39)+in_buf[158]*(-14)+in_buf[159]*(5)+in_buf[160]*(15)+in_buf[161]*(15)+in_buf[162]*(20)+in_buf[163]*(25)+in_buf[164]*(37)+in_buf[165]*(32)+in_buf[166]*(23)+in_buf[167]*(0)+in_buf[168]*(5)+in_buf[169]*(-7)+in_buf[170]*(4)+in_buf[171]*(49)+in_buf[172]*(-10)+in_buf[173]*(-12)+in_buf[174]*(4)+in_buf[175]*(-9)+in_buf[176]*(6)+in_buf[177]*(16)+in_buf[178]*(12)+in_buf[179]*(13)+in_buf[180]*(-1)+in_buf[181]*(16)+in_buf[182]*(19)+in_buf[183]*(12)+in_buf[184]*(4)+in_buf[185]*(0)+in_buf[186]*(-9)+in_buf[187]*(-9)+in_buf[188]*(17)+in_buf[189]*(17)+in_buf[190]*(-7)+in_buf[191]*(-20)+in_buf[192]*(0)+in_buf[193]*(18)+in_buf[194]*(-26)+in_buf[195]*(-8)+in_buf[196]*(1)+in_buf[197]*(-20)+in_buf[198]*(10)+in_buf[199]*(27)+in_buf[200]*(1)+in_buf[201]*(-19)+in_buf[202]*(-1)+in_buf[203]*(7)+in_buf[204]*(24)+in_buf[205]*(15)+in_buf[206]*(8)+in_buf[207]*(13)+in_buf[208]*(22)+in_buf[209]*(28)+in_buf[210]*(22)+in_buf[211]*(17)+in_buf[212]*(14)+in_buf[213]*(3)+in_buf[214]*(-2)+in_buf[215]*(5)+in_buf[216]*(14)+in_buf[217]*(0)+in_buf[218]*(-38)+in_buf[219]*(-36)+in_buf[220]*(-11)+in_buf[221]*(-10)+in_buf[222]*(-23)+in_buf[223]*(4)+in_buf[224]*(-7)+in_buf[225]*(11)+in_buf[226]*(-14)+in_buf[227]*(-20)+in_buf[228]*(-4)+in_buf[229]*(-16)+in_buf[230]*(-4)+in_buf[231]*(9)+in_buf[232]*(18)+in_buf[233]*(-1)+in_buf[234]*(19)+in_buf[235]*(22)+in_buf[236]*(16)+in_buf[237]*(14)+in_buf[238]*(30)+in_buf[239]*(19)+in_buf[240]*(26)+in_buf[241]*(6)+in_buf[242]*(2)+in_buf[243]*(-6)+in_buf[244]*(1)+in_buf[245]*(-8)+in_buf[246]*(-17)+in_buf[247]*(-46)+in_buf[248]*(-31)+in_buf[249]*(-37)+in_buf[250]*(-31)+in_buf[251]*(12)+in_buf[252]*(11)+in_buf[253]*(18)+in_buf[254]*(17)+in_buf[255]*(-14)+in_buf[256]*(-6)+in_buf[257]*(-1)+in_buf[258]*(11)+in_buf[259]*(12)+in_buf[260]*(10)+in_buf[261]*(4)+in_buf[262]*(34)+in_buf[263]*(18)+in_buf[264]*(20)+in_buf[265]*(32)+in_buf[266]*(27)+in_buf[267]*(23)+in_buf[268]*(8)+in_buf[269]*(2)+in_buf[270]*(0)+in_buf[271]*(0)+in_buf[272]*(-13)+in_buf[273]*(-8)+in_buf[274]*(-14)+in_buf[275]*(-32)+in_buf[276]*(-29)+in_buf[277]*(-39)+in_buf[278]*(-20)+in_buf[279]*(30)+in_buf[280]*(8)+in_buf[281]*(-3)+in_buf[282]*(5)+in_buf[283]*(25)+in_buf[284]*(-14)+in_buf[285]*(5)+in_buf[286]*(16)+in_buf[287]*(15)+in_buf[288]*(8)+in_buf[289]*(12)+in_buf[290]*(6)+in_buf[291]*(16)+in_buf[292]*(12)+in_buf[293]*(16)+in_buf[294]*(15)+in_buf[295]*(13)+in_buf[296]*(10)+in_buf[297]*(-9)+in_buf[298]*(0)+in_buf[299]*(3)+in_buf[300]*(-14)+in_buf[301]*(-22)+in_buf[302]*(-13)+in_buf[303]*(-20)+in_buf[304]*(-26)+in_buf[305]*(12)+in_buf[306]*(10)+in_buf[307]*(25)+in_buf[308]*(2)+in_buf[309]*(-18)+in_buf[310]*(37)+in_buf[311]*(4)+in_buf[312]*(3)+in_buf[313]*(16)+in_buf[314]*(16)+in_buf[315]*(13)+in_buf[316]*(6)+in_buf[317]*(0)+in_buf[318]*(4)+in_buf[319]*(13)+in_buf[320]*(0)+in_buf[321]*(-1)+in_buf[322]*(6)+in_buf[323]*(5)+in_buf[324]*(13)+in_buf[325]*(14)+in_buf[326]*(13)+in_buf[327]*(-11)+in_buf[328]*(-17)+in_buf[329]*(-21)+in_buf[330]*(9)+in_buf[331]*(13)+in_buf[332]*(12)+in_buf[333]*(12)+in_buf[334]*(15)+in_buf[335]*(17)+in_buf[336]*(8)+in_buf[337]*(-14)+in_buf[338]*(24)+in_buf[339]*(13)+in_buf[340]*(37)+in_buf[341]*(30)+in_buf[342]*(34)+in_buf[343]*(7)+in_buf[344]*(5)+in_buf[345]*(-2)+in_buf[346]*(-5)+in_buf[347]*(-12)+in_buf[348]*(-37)+in_buf[349]*(-20)+in_buf[350]*(1)+in_buf[351]*(5)+in_buf[352]*(5)+in_buf[353]*(18)+in_buf[354]*(3)+in_buf[355]*(-7)+in_buf[356]*(-11)+in_buf[357]*(0)+in_buf[358]*(10)+in_buf[359]*(27)+in_buf[360]*(-22)+in_buf[361]*(18)+in_buf[362]*(41)+in_buf[363]*(27)+in_buf[364]*(-18)+in_buf[365]*(-13)+in_buf[366]*(2)+in_buf[367]*(12)+in_buf[368]*(47)+in_buf[369]*(7)+in_buf[370]*(19)+in_buf[371]*(17)+in_buf[372]*(7)+in_buf[373]*(0)+in_buf[374]*(0)+in_buf[375]*(-5)+in_buf[376]*(-3)+in_buf[377]*(9)+in_buf[378]*(9)+in_buf[379]*(-6)+in_buf[380]*(3)+in_buf[381]*(1)+in_buf[382]*(-7)+in_buf[383]*(-13)+in_buf[384]*(-10)+in_buf[385]*(11)+in_buf[386]*(28)+in_buf[387]*(10)+in_buf[388]*(13)+in_buf[389]*(4)+in_buf[390]*(31)+in_buf[391]*(15)+in_buf[392]*(-13)+in_buf[393]*(-12)+in_buf[394]*(-14)+in_buf[395]*(15)+in_buf[396]*(29)+in_buf[397]*(-10)+in_buf[398]*(9)+in_buf[399]*(7)+in_buf[400]*(8)+in_buf[401]*(3)+in_buf[402]*(0)+in_buf[403]*(6)+in_buf[404]*(6)+in_buf[405]*(11)+in_buf[406]*(3)+in_buf[407]*(3)+in_buf[408]*(-5)+in_buf[409]*(-17)+in_buf[410]*(-5)+in_buf[411]*(2)+in_buf[412]*(25)+in_buf[413]*(15)+in_buf[414]*(20)+in_buf[415]*(23)+in_buf[416]*(25)+in_buf[417]*(-10)+in_buf[418]*(35)+in_buf[419]*(13)+in_buf[420]*(-15)+in_buf[421]*(-1)+in_buf[422]*(-41)+in_buf[423]*(5)+in_buf[424]*(3)+in_buf[425]*(12)+in_buf[426]*(4)+in_buf[427]*(-5)+in_buf[428]*(17)+in_buf[429]*(14)+in_buf[430]*(23)+in_buf[431]*(24)+in_buf[432]*(19)+in_buf[433]*(7)+in_buf[434]*(-3)+in_buf[435]*(0)+in_buf[436]*(-11)+in_buf[437]*(-13)+in_buf[438]*(2)+in_buf[439]*(6)+in_buf[440]*(33)+in_buf[441]*(30)+in_buf[442]*(17)+in_buf[443]*(10)+in_buf[444]*(24)+in_buf[445]*(-9)+in_buf[446]*(14)+in_buf[447]*(16)+in_buf[448]*(0)+in_buf[449]*(-1)+in_buf[450]*(-20)+in_buf[451]*(-9)+in_buf[452]*(-7)+in_buf[453]*(8)+in_buf[454]*(-2)+in_buf[455]*(0)+in_buf[456]*(13)+in_buf[457]*(7)+in_buf[458]*(16)+in_buf[459]*(33)+in_buf[460]*(21)+in_buf[461]*(8)+in_buf[462]*(-6)+in_buf[463]*(-17)+in_buf[464]*(-23)+in_buf[465]*(-5)+in_buf[466]*(3)+in_buf[467]*(14)+in_buf[468]*(24)+in_buf[469]*(22)+in_buf[470]*(22)+in_buf[471]*(12)+in_buf[472]*(1)+in_buf[473]*(-9)+in_buf[474]*(42)+in_buf[475]*(39)+in_buf[476]*(0)+in_buf[477]*(7)+in_buf[478]*(-31)+in_buf[479]*(-5)+in_buf[480]*(-25)+in_buf[481]*(0)+in_buf[482]*(-4)+in_buf[483]*(1)+in_buf[484]*(9)+in_buf[485]*(9)+in_buf[486]*(11)+in_buf[487]*(17)+in_buf[488]*(18)+in_buf[489]*(8)+in_buf[490]*(-11)+in_buf[491]*(0)+in_buf[492]*(-12)+in_buf[493]*(8)+in_buf[494]*(16)+in_buf[495]*(7)+in_buf[496]*(7)+in_buf[497]*(13)+in_buf[498]*(14)+in_buf[499]*(10)+in_buf[500]*(7)+in_buf[501]*(10)+in_buf[502]*(14)+in_buf[503]*(21)+in_buf[504]*(23)+in_buf[505]*(7)+in_buf[506]*(-20)+in_buf[507]*(-23)+in_buf[508]*(-21)+in_buf[509]*(-22)+in_buf[510]*(-11)+in_buf[511]*(-10)+in_buf[512]*(-18)+in_buf[513]*(-13)+in_buf[514]*(3)+in_buf[515]*(2)+in_buf[516]*(-13)+in_buf[517]*(-9)+in_buf[518]*(-15)+in_buf[519]*(-8)+in_buf[520]*(0)+in_buf[521]*(22)+in_buf[522]*(14)+in_buf[523]*(14)+in_buf[524]*(1)+in_buf[525]*(18)+in_buf[526]*(31)+in_buf[527]*(19)+in_buf[528]*(4)+in_buf[529]*(-1)+in_buf[530]*(28)+in_buf[531]*(-11)+in_buf[532]*(-2)+in_buf[533]*(34)+in_buf[534]*(28)+in_buf[535]*(-16)+in_buf[536]*(-22)+in_buf[537]*(-36)+in_buf[538]*(-53)+in_buf[539]*(-37)+in_buf[540]*(-31)+in_buf[541]*(-24)+in_buf[542]*(-28)+in_buf[543]*(-30)+in_buf[544]*(-16)+in_buf[545]*(-10)+in_buf[546]*(-9)+in_buf[547]*(-3)+in_buf[548]*(1)+in_buf[549]*(7)+in_buf[550]*(4)+in_buf[551]*(21)+in_buf[552]*(4)+in_buf[553]*(16)+in_buf[554]*(14)+in_buf[555]*(0)+in_buf[556]*(0)+in_buf[557]*(-4)+in_buf[558]*(4)+in_buf[559]*(-11)+in_buf[560]*(1)+in_buf[561]*(21)+in_buf[562]*(8)+in_buf[563]*(-13)+in_buf[564]*(-1)+in_buf[565]*(-36)+in_buf[566]*(-42)+in_buf[567]*(-40)+in_buf[568]*(-21)+in_buf[569]*(-34)+in_buf[570]*(-41)+in_buf[571]*(-38)+in_buf[572]*(-32)+in_buf[573]*(-6)+in_buf[574]*(-1)+in_buf[575]*(-2)+in_buf[576]*(3)+in_buf[577]*(0)+in_buf[578]*(-3)+in_buf[579]*(20)+in_buf[580]*(13)+in_buf[581]*(12)+in_buf[582]*(2)+in_buf[583]*(20)+in_buf[584]*(25)+in_buf[585]*(26)+in_buf[586]*(-5)+in_buf[587]*(-1)+in_buf[588]*(0)+in_buf[589]*(-4)+in_buf[590]*(7)+in_buf[591]*(-1)+in_buf[592]*(19)+in_buf[593]*(-28)+in_buf[594]*(-22)+in_buf[595]*(-40)+in_buf[596]*(-34)+in_buf[597]*(-38)+in_buf[598]*(-19)+in_buf[599]*(-24)+in_buf[600]*(-8)+in_buf[601]*(-12)+in_buf[602]*(-8)+in_buf[603]*(-7)+in_buf[604]*(-3)+in_buf[605]*(-13)+in_buf[606]*(10)+in_buf[607]*(-1)+in_buf[608]*(3)+in_buf[609]*(9)+in_buf[610]*(-15)+in_buf[611]*(-2)+in_buf[612]*(23)+in_buf[613]*(3)+in_buf[614]*(-14)+in_buf[615]*(0)+in_buf[616]*(2)+in_buf[617]*(-7)+in_buf[618]*(-13)+in_buf[619]*(3)+in_buf[620]*(18)+in_buf[621]*(6)+in_buf[622]*(-15)+in_buf[623]*(-47)+in_buf[624]*(-24)+in_buf[625]*(-12)+in_buf[626]*(5)+in_buf[627]*(-2)+in_buf[628]*(3)+in_buf[629]*(-9)+in_buf[630]*(-9)+in_buf[631]*(-14)+in_buf[632]*(-3)+in_buf[633]*(-12)+in_buf[634]*(-9)+in_buf[635]*(-23)+in_buf[636]*(0)+in_buf[637]*(-14)+in_buf[638]*(-5)+in_buf[639]*(15)+in_buf[640]*(35)+in_buf[641]*(11)+in_buf[642]*(2)+in_buf[643]*(1)+in_buf[644]*(4)+in_buf[645]*(0)+in_buf[646]*(-22)+in_buf[647]*(1)+in_buf[648]*(3)+in_buf[649]*(27)+in_buf[650]*(14)+in_buf[651]*(-6)+in_buf[652]*(0)+in_buf[653]*(-7)+in_buf[654]*(10)+in_buf[655]*(16)+in_buf[656]*(5)+in_buf[657]*(-8)+in_buf[658]*(-19)+in_buf[659]*(-15)+in_buf[660]*(-12)+in_buf[661]*(-13)+in_buf[662]*(-24)+in_buf[663]*(-22)+in_buf[664]*(-3)+in_buf[665]*(-18)+in_buf[666]*(2)+in_buf[667]*(13)+in_buf[668]*(51)+in_buf[669]*(16)+in_buf[670]*(-7)+in_buf[671]*(-2)+in_buf[672]*(4)+in_buf[673]*(-1)+in_buf[674]*(-2)+in_buf[675]*(1)+in_buf[676]*(19)+in_buf[677]*(34)+in_buf[678]*(16)+in_buf[679]*(13)+in_buf[680]*(33)+in_buf[681]*(23)+in_buf[682]*(26)+in_buf[683]*(6)+in_buf[684]*(-3)+in_buf[685]*(5)+in_buf[686]*(-15)+in_buf[687]*(-6)+in_buf[688]*(-6)+in_buf[689]*(6)+in_buf[690]*(-6)+in_buf[691]*(-14)+in_buf[692]*(-5)+in_buf[693]*(4)+in_buf[694]*(13)+in_buf[695]*(35)+in_buf[696]*(0)+in_buf[697]*(-11)+in_buf[698]*(-15)+in_buf[699]*(2)+in_buf[700]*(-2)+in_buf[701]*(2)+in_buf[702]*(26)+in_buf[703]*(-1)+in_buf[704]*(5)+in_buf[705]*(40)+in_buf[706]*(19)+in_buf[707]*(24)+in_buf[708]*(36)+in_buf[709]*(25)+in_buf[710]*(3)+in_buf[711]*(-3)+in_buf[712]*(9)+in_buf[713]*(8)+in_buf[714]*(-4)+in_buf[715]*(1)+in_buf[716]*(11)+in_buf[717]*(3)+in_buf[718]*(-6)+in_buf[719]*(29)+in_buf[720]*(24)+in_buf[721]*(29)+in_buf[722]*(9)+in_buf[723]*(17)+in_buf[724]*(23)+in_buf[725]*(9)+in_buf[726]*(-6)+in_buf[727]*(1)+in_buf[728]*(-2)+in_buf[729]*(3)+in_buf[730]*(0)+in_buf[731]*(9)+in_buf[732]*(10)+in_buf[733]*(39)+in_buf[734]*(52)+in_buf[735]*(44)+in_buf[736]*(23)+in_buf[737]*(35)+in_buf[738]*(53)+in_buf[739]*(27)+in_buf[740]*(39)+in_buf[741]*(63)+in_buf[742]*(84)+in_buf[743]*(40)+in_buf[744]*(52)+in_buf[745]*(41)+in_buf[746]*(37)+in_buf[747]*(55)+in_buf[748]*(67)+in_buf[749]*(49)+in_buf[750]*(53)+in_buf[751]*(10)+in_buf[752]*(21)+in_buf[753]*(-3)+in_buf[754]*(-1)+in_buf[755]*(-1)+in_buf[756]*(-3)+in_buf[757]*(-2)+in_buf[758]*(3)+in_buf[759]*(2)+in_buf[760]*(-31)+in_buf[761]*(-41)+in_buf[762]*(13)+in_buf[763]*(13)+in_buf[764]*(19)+in_buf[765]*(11)+in_buf[766]*(37)+in_buf[767]*(31)+in_buf[768]*(29)+in_buf[769]*(1)+in_buf[770]*(47)+in_buf[771]*(36)+in_buf[772]*(27)+in_buf[773]*(5)+in_buf[774]*(16)+in_buf[775]*(39)+in_buf[776]*(22)+in_buf[777]*(23)+in_buf[778]*(25)+in_buf[779]*(-3)+in_buf[780]*(-3)+in_buf[781]*(2)+in_buf[782]*(0)+in_buf[783]*(-2);
assign in_buf_weight038=in_buf[0]*(1)+in_buf[1]*(0)+in_buf[2]*(4)+in_buf[3]*(-3)+in_buf[4]*(4)+in_buf[5]*(2)+in_buf[6]*(3)+in_buf[7]*(3)+in_buf[8]*(3)+in_buf[9]*(5)+in_buf[10]*(-3)+in_buf[11]*(0)+in_buf[12]*(-11)+in_buf[13]*(-6)+in_buf[14]*(5)+in_buf[15]*(10)+in_buf[16]*(3)+in_buf[17]*(3)+in_buf[18]*(2)+in_buf[19]*(4)+in_buf[20]*(3)+in_buf[21]*(-2)+in_buf[22]*(0)+in_buf[23]*(1)+in_buf[24]*(3)+in_buf[25]*(0)+in_buf[26]*(-3)+in_buf[27]*(3)+in_buf[28]*(-2)+in_buf[29]*(0)+in_buf[30]*(3)+in_buf[31]*(0)+in_buf[32]*(-5)+in_buf[33]*(1)+in_buf[34]*(-1)+in_buf[35]*(-2)+in_buf[36]*(-7)+in_buf[37]*(-7)+in_buf[38]*(-3)+in_buf[39]*(10)+in_buf[40]*(-1)+in_buf[41]*(-20)+in_buf[42]*(-4)+in_buf[43]*(-9)+in_buf[44]*(19)+in_buf[45]*(-5)+in_buf[46]*(-21)+in_buf[47]*(-21)+in_buf[48]*(-27)+in_buf[49]*(-27)+in_buf[50]*(-15)+in_buf[51]*(-11)+in_buf[52]*(1)+in_buf[53]*(4)+in_buf[54]*(1)+in_buf[55]*(2)+in_buf[56]*(0)+in_buf[57]*(4)+in_buf[58]*(-18)+in_buf[59]*(4)+in_buf[60]*(-12)+in_buf[61]*(-1)+in_buf[62]*(-17)+in_buf[63]*(-10)+in_buf[64]*(13)+in_buf[65]*(31)+in_buf[66]*(31)+in_buf[67]*(7)+in_buf[68]*(9)+in_buf[69]*(-8)+in_buf[70]*(-4)+in_buf[71]*(-15)+in_buf[72]*(-21)+in_buf[73]*(-32)+in_buf[74]*(-24)+in_buf[75]*(-34)+in_buf[76]*(-9)+in_buf[77]*(0)+in_buf[78]*(-23)+in_buf[79]*(-6)+in_buf[80]*(10)+in_buf[81]*(8)+in_buf[82]*(-3)+in_buf[83]*(-4)+in_buf[84]*(-4)+in_buf[85]*(1)+in_buf[86]*(-20)+in_buf[87]*(1)+in_buf[88]*(-20)+in_buf[89]*(8)+in_buf[90]*(-4)+in_buf[91]*(-10)+in_buf[92]*(-1)+in_buf[93]*(15)+in_buf[94]*(7)+in_buf[95]*(24)+in_buf[96]*(9)+in_buf[97]*(12)+in_buf[98]*(8)+in_buf[99]*(10)+in_buf[100]*(8)+in_buf[101]*(-6)+in_buf[102]*(-10)+in_buf[103]*(-20)+in_buf[104]*(-37)+in_buf[105]*(-22)+in_buf[106]*(-23)+in_buf[107]*(-5)+in_buf[108]*(-2)+in_buf[109]*(-8)+in_buf[110]*(-22)+in_buf[111]*(-2)+in_buf[112]*(3)+in_buf[113]*(-1)+in_buf[114]*(-25)+in_buf[115]*(-37)+in_buf[116]*(-30)+in_buf[117]*(-14)+in_buf[118]*(1)+in_buf[119]*(11)+in_buf[120]*(14)+in_buf[121]*(16)+in_buf[122]*(11)+in_buf[123]*(13)+in_buf[124]*(17)+in_buf[125]*(0)+in_buf[126]*(5)+in_buf[127]*(-2)+in_buf[128]*(11)+in_buf[129]*(19)+in_buf[130]*(-3)+in_buf[131]*(-20)+in_buf[132]*(-14)+in_buf[133]*(-26)+in_buf[134]*(-30)+in_buf[135]*(-33)+in_buf[136]*(-10)+in_buf[137]*(15)+in_buf[138]*(22)+in_buf[139]*(3)+in_buf[140]*(0)+in_buf[141]*(1)+in_buf[142]*(-27)+in_buf[143]*(-4)+in_buf[144]*(-7)+in_buf[145]*(-45)+in_buf[146]*(-25)+in_buf[147]*(-4)+in_buf[148]*(-12)+in_buf[149]*(-1)+in_buf[150]*(10)+in_buf[151]*(21)+in_buf[152]*(20)+in_buf[153]*(-1)+in_buf[154]*(5)+in_buf[155]*(7)+in_buf[156]*(16)+in_buf[157]*(25)+in_buf[158]*(13)+in_buf[159]*(14)+in_buf[160]*(14)+in_buf[161]*(-1)+in_buf[162]*(-10)+in_buf[163]*(-21)+in_buf[164]*(-10)+in_buf[165]*(17)+in_buf[166]*(16)+in_buf[167]*(-13)+in_buf[168]*(0)+in_buf[169]*(10)+in_buf[170]*(11)+in_buf[171]*(-19)+in_buf[172]*(-8)+in_buf[173]*(-38)+in_buf[174]*(-29)+in_buf[175]*(-7)+in_buf[176]*(-16)+in_buf[177]*(-5)+in_buf[178]*(6)+in_buf[179]*(2)+in_buf[180]*(0)+in_buf[181]*(-7)+in_buf[182]*(-10)+in_buf[183]*(-8)+in_buf[184]*(6)+in_buf[185]*(8)+in_buf[186]*(3)+in_buf[187]*(-5)+in_buf[188]*(-4)+in_buf[189]*(-4)+in_buf[190]*(-5)+in_buf[191]*(-4)+in_buf[192]*(-28)+in_buf[193]*(-6)+in_buf[194]*(-12)+in_buf[195]*(-30)+in_buf[196]*(-9)+in_buf[197]*(-15)+in_buf[198]*(11)+in_buf[199]*(-30)+in_buf[200]*(17)+in_buf[201]*(2)+in_buf[202]*(0)+in_buf[203]*(-1)+in_buf[204]*(18)+in_buf[205]*(-2)+in_buf[206]*(-3)+in_buf[207]*(-1)+in_buf[208]*(-18)+in_buf[209]*(-14)+in_buf[210]*(-15)+in_buf[211]*(0)+in_buf[212]*(-2)+in_buf[213]*(-7)+in_buf[214]*(2)+in_buf[215]*(3)+in_buf[216]*(-17)+in_buf[217]*(7)+in_buf[218]*(14)+in_buf[219]*(-2)+in_buf[220]*(-5)+in_buf[221]*(11)+in_buf[222]*(-21)+in_buf[223]*(-34)+in_buf[224]*(24)+in_buf[225]*(-22)+in_buf[226]*(15)+in_buf[227]*(17)+in_buf[228]*(26)+in_buf[229]*(4)+in_buf[230]*(1)+in_buf[231]*(-8)+in_buf[232]*(0)+in_buf[233]*(-7)+in_buf[234]*(-8)+in_buf[235]*(-13)+in_buf[236]*(-11)+in_buf[237]*(7)+in_buf[238]*(4)+in_buf[239]*(0)+in_buf[240]*(4)+in_buf[241]*(1)+in_buf[242]*(2)+in_buf[243]*(7)+in_buf[244]*(-3)+in_buf[245]*(10)+in_buf[246]*(8)+in_buf[247]*(3)+in_buf[248]*(1)+in_buf[249]*(4)+in_buf[250]*(3)+in_buf[251]*(13)+in_buf[252]*(-8)+in_buf[253]*(-30)+in_buf[254]*(15)+in_buf[255]*(39)+in_buf[256]*(16)+in_buf[257]*(2)+in_buf[258]*(5)+in_buf[259]*(-13)+in_buf[260]*(-16)+in_buf[261]*(0)+in_buf[262]*(-4)+in_buf[263]*(-13)+in_buf[264]*(-2)+in_buf[265]*(12)+in_buf[266]*(11)+in_buf[267]*(4)+in_buf[268]*(3)+in_buf[269]*(-3)+in_buf[270]*(-6)+in_buf[271]*(0)+in_buf[272]*(0)+in_buf[273]*(-2)+in_buf[274]*(1)+in_buf[275]*(5)+in_buf[276]*(-8)+in_buf[277]*(-9)+in_buf[278]*(-10)+in_buf[279]*(-25)+in_buf[280]*(-10)+in_buf[281]*(-28)+in_buf[282]*(12)+in_buf[283]*(55)+in_buf[284]*(19)+in_buf[285]*(24)+in_buf[286]*(17)+in_buf[287]*(-9)+in_buf[288]*(-20)+in_buf[289]*(-2)+in_buf[290]*(0)+in_buf[291]*(3)+in_buf[292]*(11)+in_buf[293]*(-5)+in_buf[294]*(-2)+in_buf[295]*(-11)+in_buf[296]*(-14)+in_buf[297]*(-11)+in_buf[298]*(-8)+in_buf[299]*(-11)+in_buf[300]*(-3)+in_buf[301]*(3)+in_buf[302]*(12)+in_buf[303]*(32)+in_buf[304]*(-13)+in_buf[305]*(-49)+in_buf[306]*(-12)+in_buf[307]*(-8)+in_buf[308]*(-20)+in_buf[309]*(-7)+in_buf[310]*(18)+in_buf[311]*(36)+in_buf[312]*(19)+in_buf[313]*(17)+in_buf[314]*(13)+in_buf[315]*(-5)+in_buf[316]*(-18)+in_buf[317]*(-3)+in_buf[318]*(0)+in_buf[319]*(4)+in_buf[320]*(-3)+in_buf[321]*(-20)+in_buf[322]*(-18)+in_buf[323]*(-28)+in_buf[324]*(-15)+in_buf[325]*(-14)+in_buf[326]*(-21)+in_buf[327]*(1)+in_buf[328]*(4)+in_buf[329]*(25)+in_buf[330]*(25)+in_buf[331]*(28)+in_buf[332]*(24)+in_buf[333]*(9)+in_buf[334]*(14)+in_buf[335]*(-30)+in_buf[336]*(-19)+in_buf[337]*(-9)+in_buf[338]*(24)+in_buf[339]*(10)+in_buf[340]*(20)+in_buf[341]*(8)+in_buf[342]*(2)+in_buf[343]*(-20)+in_buf[344]*(-20)+in_buf[345]*(-2)+in_buf[346]*(-17)+in_buf[347]*(-16)+in_buf[348]*(-16)+in_buf[349]*(-29)+in_buf[350]*(-30)+in_buf[351]*(-21)+in_buf[352]*(-10)+in_buf[353]*(-8)+in_buf[354]*(-14)+in_buf[355]*(6)+in_buf[356]*(12)+in_buf[357]*(20)+in_buf[358]*(3)+in_buf[359]*(34)+in_buf[360]*(48)+in_buf[361]*(18)+in_buf[362]*(-3)+in_buf[363]*(-29)+in_buf[364]*(5)+in_buf[365]*(13)+in_buf[366]*(0)+in_buf[367]*(-4)+in_buf[368]*(0)+in_buf[369]*(-6)+in_buf[370]*(-9)+in_buf[371]*(-5)+in_buf[372]*(2)+in_buf[373]*(2)+in_buf[374]*(2)+in_buf[375]*(-6)+in_buf[376]*(0)+in_buf[377]*(-8)+in_buf[378]*(-11)+in_buf[379]*(1)+in_buf[380]*(-2)+in_buf[381]*(-6)+in_buf[382]*(2)+in_buf[383]*(10)+in_buf[384]*(13)+in_buf[385]*(6)+in_buf[386]*(26)+in_buf[387]*(42)+in_buf[388]*(25)+in_buf[389]*(39)+in_buf[390]*(39)+in_buf[391]*(22)+in_buf[392]*(-10)+in_buf[393]*(0)+in_buf[394]*(-6)+in_buf[395]*(-6)+in_buf[396]*(1)+in_buf[397]*(-5)+in_buf[398]*(3)+in_buf[399]*(-2)+in_buf[400]*(-2)+in_buf[401]*(2)+in_buf[402]*(7)+in_buf[403]*(17)+in_buf[404]*(12)+in_buf[405]*(10)+in_buf[406]*(7)+in_buf[407]*(4)+in_buf[408]*(9)+in_buf[409]*(0)+in_buf[410]*(5)+in_buf[411]*(5)+in_buf[412]*(3)+in_buf[413]*(15)+in_buf[414]*(18)+in_buf[415]*(2)+in_buf[416]*(11)+in_buf[417]*(56)+in_buf[418]*(56)+in_buf[419]*(19)+in_buf[420]*(-6)+in_buf[421]*(-5)+in_buf[422]*(-8)+in_buf[423]*(20)+in_buf[424]*(8)+in_buf[425]*(6)+in_buf[426]*(-9)+in_buf[427]*(-1)+in_buf[428]*(11)+in_buf[429]*(17)+in_buf[430]*(15)+in_buf[431]*(17)+in_buf[432]*(14)+in_buf[433]*(21)+in_buf[434]*(15)+in_buf[435]*(13)+in_buf[436]*(19)+in_buf[437]*(1)+in_buf[438]*(2)+in_buf[439]*(6)+in_buf[440]*(-4)+in_buf[441]*(-13)+in_buf[442]*(-5)+in_buf[443]*(-3)+in_buf[444]*(23)+in_buf[445]*(36)+in_buf[446]*(19)+in_buf[447]*(30)+in_buf[448]*(5)+in_buf[449]*(-2)+in_buf[450]*(-4)+in_buf[451]*(20)+in_buf[452]*(-5)+in_buf[453]*(7)+in_buf[454]*(9)+in_buf[455]*(0)+in_buf[456]*(10)+in_buf[457]*(14)+in_buf[458]*(29)+in_buf[459]*(24)+in_buf[460]*(19)+in_buf[461]*(11)+in_buf[462]*(15)+in_buf[463]*(14)+in_buf[464]*(11)+in_buf[465]*(13)+in_buf[466]*(6)+in_buf[467]*(5)+in_buf[468]*(-9)+in_buf[469]*(2)+in_buf[470]*(10)+in_buf[471]*(9)+in_buf[472]*(2)+in_buf[473]*(37)+in_buf[474]*(59)+in_buf[475]*(36)+in_buf[476]*(3)+in_buf[477]*(-6)+in_buf[478]*(4)+in_buf[479]*(12)+in_buf[480]*(6)+in_buf[481]*(1)+in_buf[482]*(10)+in_buf[483]*(3)+in_buf[484]*(10)+in_buf[485]*(15)+in_buf[486]*(21)+in_buf[487]*(15)+in_buf[488]*(25)+in_buf[489]*(18)+in_buf[490]*(11)+in_buf[491]*(12)+in_buf[492]*(8)+in_buf[493]*(11)+in_buf[494]*(-7)+in_buf[495]*(-7)+in_buf[496]*(-5)+in_buf[497]*(-1)+in_buf[498]*(1)+in_buf[499]*(0)+in_buf[500]*(5)+in_buf[501]*(18)+in_buf[502]*(31)+in_buf[503]*(48)+in_buf[504]*(3)+in_buf[505]*(-7)+in_buf[506]*(5)+in_buf[507]*(2)+in_buf[508]*(13)+in_buf[509]*(7)+in_buf[510]*(12)+in_buf[511]*(24)+in_buf[512]*(5)+in_buf[513]*(7)+in_buf[514]*(15)+in_buf[515]*(6)+in_buf[516]*(18)+in_buf[517]*(15)+in_buf[518]*(16)+in_buf[519]*(4)+in_buf[520]*(0)+in_buf[521]*(2)+in_buf[522]*(-1)+in_buf[523]*(1)+in_buf[524]*(3)+in_buf[525]*(-8)+in_buf[526]*(7)+in_buf[527]*(14)+in_buf[528]*(14)+in_buf[529]*(23)+in_buf[530]*(8)+in_buf[531]*(32)+in_buf[532]*(-4)+in_buf[533]*(-2)+in_buf[534]*(-3)+in_buf[535]*(-1)+in_buf[536]*(20)+in_buf[537]*(26)+in_buf[538]*(9)+in_buf[539]*(19)+in_buf[540]*(8)+in_buf[541]*(6)+in_buf[542]*(22)+in_buf[543]*(10)+in_buf[544]*(10)+in_buf[545]*(17)+in_buf[546]*(9)+in_buf[547]*(9)+in_buf[548]*(3)+in_buf[549]*(9)+in_buf[550]*(7)+in_buf[551]*(10)+in_buf[552]*(-4)+in_buf[553]*(-1)+in_buf[554]*(26)+in_buf[555]*(32)+in_buf[556]*(13)+in_buf[557]*(15)+in_buf[558]*(63)+in_buf[559]*(11)+in_buf[560]*(3)+in_buf[561]*(-1)+in_buf[562]*(15)+in_buf[563]*(19)+in_buf[564]*(23)+in_buf[565]*(30)+in_buf[566]*(16)+in_buf[567]*(24)+in_buf[568]*(9)+in_buf[569]*(0)+in_buf[570]*(11)+in_buf[571]*(14)+in_buf[572]*(10)+in_buf[573]*(6)+in_buf[574]*(0)+in_buf[575]*(10)+in_buf[576]*(-12)+in_buf[577]*(-7)+in_buf[578]*(8)+in_buf[579]*(-4)+in_buf[580]*(8)+in_buf[581]*(18)+in_buf[582]*(6)+in_buf[583]*(23)+in_buf[584]*(8)+in_buf[585]*(32)+in_buf[586]*(39)+in_buf[587]*(-2)+in_buf[588]*(-17)+in_buf[589]*(10)+in_buf[590]*(27)+in_buf[591]*(30)+in_buf[592]*(38)+in_buf[593]*(15)+in_buf[594]*(21)+in_buf[595]*(15)+in_buf[596]*(5)+in_buf[597]*(7)+in_buf[598]*(3)+in_buf[599]*(6)+in_buf[600]*(1)+in_buf[601]*(8)+in_buf[602]*(0)+in_buf[603]*(0)+in_buf[604]*(1)+in_buf[605]*(11)+in_buf[606]*(0)+in_buf[607]*(1)+in_buf[608]*(-4)+in_buf[609]*(-2)+in_buf[610]*(29)+in_buf[611]*(36)+in_buf[612]*(-4)+in_buf[613]*(8)+in_buf[614]*(35)+in_buf[615]*(3)+in_buf[616]*(-18)+in_buf[617]*(-11)+in_buf[618]*(21)+in_buf[619]*(12)+in_buf[620]*(27)+in_buf[621]*(9)+in_buf[622]*(17)+in_buf[623]*(15)+in_buf[624]*(6)+in_buf[625]*(5)+in_buf[626]*(-1)+in_buf[627]*(15)+in_buf[628]*(10)+in_buf[629]*(10)+in_buf[630]*(2)+in_buf[631]*(-10)+in_buf[632]*(-4)+in_buf[633]*(6)+in_buf[634]*(5)+in_buf[635]*(6)+in_buf[636]*(0)+in_buf[637]*(5)+in_buf[638]*(28)+in_buf[639]*(33)+in_buf[640]*(33)+in_buf[641]*(11)+in_buf[642]*(-26)+in_buf[643]*(5)+in_buf[644]*(4)+in_buf[645]*(0)+in_buf[646]*(18)+in_buf[647]*(17)+in_buf[648]*(4)+in_buf[649]*(-4)+in_buf[650]*(3)+in_buf[651]*(0)+in_buf[652]*(12)+in_buf[653]*(-4)+in_buf[654]*(-4)+in_buf[655]*(7)+in_buf[656]*(-2)+in_buf[657]*(4)+in_buf[658]*(0)+in_buf[659]*(5)+in_buf[660]*(5)+in_buf[661]*(8)+in_buf[662]*(19)+in_buf[663]*(6)+in_buf[664]*(18)+in_buf[665]*(27)+in_buf[666]*(40)+in_buf[667]*(41)+in_buf[668]*(19)+in_buf[669]*(1)+in_buf[670]*(-31)+in_buf[671]*(-3)+in_buf[672]*(4)+in_buf[673]*(2)+in_buf[674]*(-3)+in_buf[675]*(-2)+in_buf[676]*(-12)+in_buf[677]*(-21)+in_buf[678]*(-6)+in_buf[679]*(-9)+in_buf[680]*(-3)+in_buf[681]*(-6)+in_buf[682]*(-18)+in_buf[683]*(-5)+in_buf[684]*(11)+in_buf[685]*(3)+in_buf[686]*(1)+in_buf[687]*(2)+in_buf[688]*(11)+in_buf[689]*(-7)+in_buf[690]*(3)+in_buf[691]*(17)+in_buf[692]*(22)+in_buf[693]*(4)+in_buf[694]*(22)+in_buf[695]*(39)+in_buf[696]*(27)+in_buf[697]*(13)+in_buf[698]*(3)+in_buf[699]*(-1)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(16)+in_buf[703]*(-28)+in_buf[704]*(-26)+in_buf[705]*(-18)+in_buf[706]*(-3)+in_buf[707]*(7)+in_buf[708]*(-3)+in_buf[709]*(-16)+in_buf[710]*(-16)+in_buf[711]*(-19)+in_buf[712]*(-29)+in_buf[713]*(0)+in_buf[714]*(8)+in_buf[715]*(4)+in_buf[716]*(0)+in_buf[717]*(-9)+in_buf[718]*(0)+in_buf[719]*(18)+in_buf[720]*(2)+in_buf[721]*(-21)+in_buf[722]*(-24)+in_buf[723]*(-17)+in_buf[724]*(-22)+in_buf[725]*(0)+in_buf[726]*(7)+in_buf[727]*(-2)+in_buf[728]*(1)+in_buf[729]*(-3)+in_buf[730]*(1)+in_buf[731]*(-2)+in_buf[732]*(35)+in_buf[733]*(28)+in_buf[734]*(16)+in_buf[735]*(5)+in_buf[736]*(11)+in_buf[737]*(-15)+in_buf[738]*(-17)+in_buf[739]*(4)+in_buf[740]*(17)+in_buf[741]*(10)+in_buf[742]*(2)+in_buf[743]*(-4)+in_buf[744]*(3)+in_buf[745]*(-15)+in_buf[746]*(7)+in_buf[747]*(19)+in_buf[748]*(1)+in_buf[749]*(-15)+in_buf[750]*(4)+in_buf[751]*(18)+in_buf[752]*(42)+in_buf[753]*(-12)+in_buf[754]*(4)+in_buf[755]*(3)+in_buf[756]*(-4)+in_buf[757]*(4)+in_buf[758]*(-3)+in_buf[759]*(0)+in_buf[760]*(-29)+in_buf[761]*(-12)+in_buf[762]*(-2)+in_buf[763]*(11)+in_buf[764]*(13)+in_buf[765]*(6)+in_buf[766]*(21)+in_buf[767]*(21)+in_buf[768]*(21)+in_buf[769]*(0)+in_buf[770]*(3)+in_buf[771]*(-10)+in_buf[772]*(-5)+in_buf[773]*(-10)+in_buf[774]*(-9)+in_buf[775]*(27)+in_buf[776]*(5)+in_buf[777]*(-8)+in_buf[778]*(-19)+in_buf[779]*(-23)+in_buf[780]*(-2)+in_buf[781]*(1)+in_buf[782]*(2)+in_buf[783]*(3);
assign in_buf_weight039=in_buf[0]*(0)+in_buf[1]*(4)+in_buf[2]*(-1)+in_buf[3]*(3)+in_buf[4]*(-1)+in_buf[5]*(4)+in_buf[6]*(1)+in_buf[7]*(4)+in_buf[8]*(0)+in_buf[9]*(0)+in_buf[10]*(2)+in_buf[11]*(0)+in_buf[12]*(16)+in_buf[13]*(7)+in_buf[14]*(-17)+in_buf[15]*(-14)+in_buf[16]*(0)+in_buf[17]*(4)+in_buf[18]*(2)+in_buf[19]*(4)+in_buf[20]*(-2)+in_buf[21]*(0)+in_buf[22]*(-3)+in_buf[23]*(-2)+in_buf[24]*(3)+in_buf[25]*(0)+in_buf[26]*(4)+in_buf[27]*(4)+in_buf[28]*(1)+in_buf[29]*(-1)+in_buf[30]*(5)+in_buf[31]*(0)+in_buf[32]*(5)+in_buf[33]*(-4)+in_buf[34]*(-1)+in_buf[35]*(4)+in_buf[36]*(8)+in_buf[37]*(13)+in_buf[38]*(17)+in_buf[39]*(20)+in_buf[40]*(21)+in_buf[41]*(26)+in_buf[42]*(6)+in_buf[43]*(21)+in_buf[44]*(20)+in_buf[45]*(32)+in_buf[46]*(17)+in_buf[47]*(12)+in_buf[48]*(20)+in_buf[49]*(13)+in_buf[50]*(16)+in_buf[51]*(6)+in_buf[52]*(-3)+in_buf[53]*(-1)+in_buf[54]*(-3)+in_buf[55]*(0)+in_buf[56]*(-2)+in_buf[57]*(3)+in_buf[58]*(14)+in_buf[59]*(29)+in_buf[60]*(29)+in_buf[61]*(-6)+in_buf[62]*(0)+in_buf[63]*(13)+in_buf[64]*(-12)+in_buf[65]*(-36)+in_buf[66]*(-38)+in_buf[67]*(-13)+in_buf[68]*(-33)+in_buf[69]*(-50)+in_buf[70]*(-38)+in_buf[71]*(-29)+in_buf[72]*(-21)+in_buf[73]*(-5)+in_buf[74]*(5)+in_buf[75]*(-22)+in_buf[76]*(-25)+in_buf[77]*(-21)+in_buf[78]*(-7)+in_buf[79]*(-27)+in_buf[80]*(-13)+in_buf[81]*(-12)+in_buf[82]*(1)+in_buf[83]*(3)+in_buf[84]*(0)+in_buf[85]*(-3)+in_buf[86]*(-19)+in_buf[87]*(22)+in_buf[88]*(22)+in_buf[89]*(-5)+in_buf[90]*(-18)+in_buf[91]*(-24)+in_buf[92]*(-40)+in_buf[93]*(-27)+in_buf[94]*(-24)+in_buf[95]*(-45)+in_buf[96]*(-45)+in_buf[97]*(-11)+in_buf[98]*(9)+in_buf[99]*(1)+in_buf[100]*(-13)+in_buf[101]*(-2)+in_buf[102]*(-8)+in_buf[103]*(-29)+in_buf[104]*(1)+in_buf[105]*(9)+in_buf[106]*(0)+in_buf[107]*(42)+in_buf[108]*(11)+in_buf[109]*(-7)+in_buf[110]*(11)+in_buf[111]*(1)+in_buf[112]*(2)+in_buf[113]*(-3)+in_buf[114]*(-23)+in_buf[115]*(5)+in_buf[116]*(0)+in_buf[117]*(-53)+in_buf[118]*(-50)+in_buf[119]*(-12)+in_buf[120]*(-34)+in_buf[121]*(-17)+in_buf[122]*(-12)+in_buf[123]*(-12)+in_buf[124]*(-6)+in_buf[125]*(-6)+in_buf[126]*(9)+in_buf[127]*(6)+in_buf[128]*(7)+in_buf[129]*(7)+in_buf[130]*(-5)+in_buf[131]*(-12)+in_buf[132]*(-7)+in_buf[133]*(8)+in_buf[134]*(-3)+in_buf[135]*(24)+in_buf[136]*(38)+in_buf[137]*(27)+in_buf[138]*(37)+in_buf[139]*(28)+in_buf[140]*(0)+in_buf[141]*(2)+in_buf[142]*(-5)+in_buf[143]*(-30)+in_buf[144]*(-26)+in_buf[145]*(-38)+in_buf[146]*(-14)+in_buf[147]*(-4)+in_buf[148]*(-4)+in_buf[149]*(9)+in_buf[150]*(17)+in_buf[151]*(22)+in_buf[152]*(18)+in_buf[153]*(22)+in_buf[154]*(22)+in_buf[155]*(4)+in_buf[156]*(10)+in_buf[157]*(22)+in_buf[158]*(3)+in_buf[159]*(3)+in_buf[160]*(5)+in_buf[161]*(10)+in_buf[162]*(-4)+in_buf[163]*(-13)+in_buf[164]*(-7)+in_buf[165]*(21)+in_buf[166]*(47)+in_buf[167]*(26)+in_buf[168]*(-3)+in_buf[169]*(-22)+in_buf[170]*(4)+in_buf[171]*(-56)+in_buf[172]*(-37)+in_buf[173]*(0)+in_buf[174]*(-13)+in_buf[175]*(1)+in_buf[176]*(6)+in_buf[177]*(-1)+in_buf[178]*(6)+in_buf[179]*(15)+in_buf[180]*(12)+in_buf[181]*(16)+in_buf[182]*(17)+in_buf[183]*(10)+in_buf[184]*(9)+in_buf[185]*(20)+in_buf[186]*(6)+in_buf[187]*(12)+in_buf[188]*(5)+in_buf[189]*(8)+in_buf[190]*(16)+in_buf[191]*(17)+in_buf[192]*(21)+in_buf[193]*(26)+in_buf[194]*(-1)+in_buf[195]*(-14)+in_buf[196]*(1)+in_buf[197]*(-45)+in_buf[198]*(0)+in_buf[199]*(-62)+in_buf[200]*(-36)+in_buf[201]*(12)+in_buf[202]*(-3)+in_buf[203]*(-15)+in_buf[204]*(11)+in_buf[205]*(17)+in_buf[206]*(19)+in_buf[207]*(15)+in_buf[208]*(4)+in_buf[209]*(-2)+in_buf[210]*(-2)+in_buf[211]*(16)+in_buf[212]*(12)+in_buf[213]*(8)+in_buf[214]*(13)+in_buf[215]*(5)+in_buf[216]*(-5)+in_buf[217]*(6)+in_buf[218]*(19)+in_buf[219]*(24)+in_buf[220]*(20)+in_buf[221]*(42)+in_buf[222]*(-2)+in_buf[223]*(-16)+in_buf[224]*(26)+in_buf[225]*(-42)+in_buf[226]*(-8)+in_buf[227]*(-4)+in_buf[228]*(-15)+in_buf[229]*(3)+in_buf[230]*(16)+in_buf[231]*(3)+in_buf[232]*(24)+in_buf[233]*(21)+in_buf[234]*(8)+in_buf[235]*(11)+in_buf[236]*(7)+in_buf[237]*(9)+in_buf[238]*(1)+in_buf[239]*(2)+in_buf[240]*(21)+in_buf[241]*(7)+in_buf[242]*(12)+in_buf[243]*(7)+in_buf[244]*(6)+in_buf[245]*(10)+in_buf[246]*(2)+in_buf[247]*(0)+in_buf[248]*(41)+in_buf[249]*(41)+in_buf[250]*(3)+in_buf[251]*(17)+in_buf[252]*(-6)+in_buf[253]*(-9)+in_buf[254]*(-7)+in_buf[255]*(2)+in_buf[256]*(-18)+in_buf[257]*(-5)+in_buf[258]*(18)+in_buf[259]*(8)+in_buf[260]*(9)+in_buf[261]*(19)+in_buf[262]*(11)+in_buf[263]*(12)+in_buf[264]*(-1)+in_buf[265]*(14)+in_buf[266]*(3)+in_buf[267]*(-13)+in_buf[268]*(-1)+in_buf[269]*(4)+in_buf[270]*(0)+in_buf[271]*(1)+in_buf[272]*(4)+in_buf[273]*(2)+in_buf[274]*(-17)+in_buf[275]*(2)+in_buf[276]*(37)+in_buf[277]*(60)+in_buf[278]*(-2)+in_buf[279]*(-18)+in_buf[280]*(-6)+in_buf[281]*(-8)+in_buf[282]*(-2)+in_buf[283]*(-4)+in_buf[284]*(10)+in_buf[285]*(4)+in_buf[286]*(14)+in_buf[287]*(20)+in_buf[288]*(17)+in_buf[289]*(17)+in_buf[290]*(13)+in_buf[291]*(6)+in_buf[292]*(15)+in_buf[293]*(11)+in_buf[294]*(7)+in_buf[295]*(-2)+in_buf[296]*(-6)+in_buf[297]*(-4)+in_buf[298]*(0)+in_buf[299]*(-12)+in_buf[300]*(0)+in_buf[301]*(0)+in_buf[302]*(1)+in_buf[303]*(15)+in_buf[304]*(29)+in_buf[305]*(10)+in_buf[306]*(17)+in_buf[307]*(-7)+in_buf[308]*(-9)+in_buf[309]*(9)+in_buf[310]*(-38)+in_buf[311]*(-2)+in_buf[312]*(3)+in_buf[313]*(2)+in_buf[314]*(30)+in_buf[315]*(21)+in_buf[316]*(17)+in_buf[317]*(12)+in_buf[318]*(13)+in_buf[319]*(10)+in_buf[320]*(15)+in_buf[321]*(15)+in_buf[322]*(9)+in_buf[323]*(0)+in_buf[324]*(-4)+in_buf[325]*(0)+in_buf[326]*(-6)+in_buf[327]*(-14)+in_buf[328]*(-7)+in_buf[329]*(16)+in_buf[330]*(-4)+in_buf[331]*(7)+in_buf[332]*(25)+in_buf[333]*(16)+in_buf[334]*(59)+in_buf[335]*(-18)+in_buf[336]*(-10)+in_buf[337]*(-14)+in_buf[338]*(-10)+in_buf[339]*(14)+in_buf[340]*(8)+in_buf[341]*(9)+in_buf[342]*(30)+in_buf[343]*(20)+in_buf[344]*(4)+in_buf[345]*(15)+in_buf[346]*(8)+in_buf[347]*(8)+in_buf[348]*(9)+in_buf[349]*(13)+in_buf[350]*(-13)+in_buf[351]*(-7)+in_buf[352]*(-10)+in_buf[353]*(1)+in_buf[354]*(-10)+in_buf[355]*(11)+in_buf[356]*(12)+in_buf[357]*(19)+in_buf[358]*(0)+in_buf[359]*(16)+in_buf[360]*(19)+in_buf[361]*(-4)+in_buf[362]*(15)+in_buf[363]*(-36)+in_buf[364]*(-13)+in_buf[365]*(-4)+in_buf[366]*(-19)+in_buf[367]*(22)+in_buf[368]*(12)+in_buf[369]*(8)+in_buf[370]*(16)+in_buf[371]*(26)+in_buf[372]*(5)+in_buf[373]*(18)+in_buf[374]*(9)+in_buf[375]*(20)+in_buf[376]*(15)+in_buf[377]*(1)+in_buf[378]*(0)+in_buf[379]*(5)+in_buf[380]*(-6)+in_buf[381]*(-11)+in_buf[382]*(6)+in_buf[383]*(23)+in_buf[384]*(14)+in_buf[385]*(5)+in_buf[386]*(12)+in_buf[387]*(30)+in_buf[388]*(-8)+in_buf[389]*(2)+in_buf[390]*(0)+in_buf[391]*(-8)+in_buf[392]*(14)+in_buf[393]*(-10)+in_buf[394]*(-28)+in_buf[395]*(2)+in_buf[396]*(-1)+in_buf[397]*(13)+in_buf[398]*(15)+in_buf[399]*(7)+in_buf[400]*(8)+in_buf[401]*(11)+in_buf[402]*(9)+in_buf[403]*(25)+in_buf[404]*(13)+in_buf[405]*(9)+in_buf[406]*(-6)+in_buf[407]*(0)+in_buf[408]*(-14)+in_buf[409]*(-5)+in_buf[410]*(0)+in_buf[411]*(4)+in_buf[412]*(8)+in_buf[413]*(7)+in_buf[414]*(1)+in_buf[415]*(20)+in_buf[416]*(17)+in_buf[417]*(8)+in_buf[418]*(-35)+in_buf[419]*(-22)+in_buf[420]*(8)+in_buf[421]*(-14)+in_buf[422]*(-13)+in_buf[423]*(-18)+in_buf[424]*(-4)+in_buf[425]*(-11)+in_buf[426]*(0)+in_buf[427]*(19)+in_buf[428]*(17)+in_buf[429]*(15)+in_buf[430]*(15)+in_buf[431]*(17)+in_buf[432]*(7)+in_buf[433]*(-3)+in_buf[434]*(-5)+in_buf[435]*(-10)+in_buf[436]*(-4)+in_buf[437]*(-6)+in_buf[438]*(-6)+in_buf[439]*(-7)+in_buf[440]*(5)+in_buf[441]*(-2)+in_buf[442]*(6)+in_buf[443]*(18)+in_buf[444]*(17)+in_buf[445]*(25)+in_buf[446]*(-16)+in_buf[447]*(-21)+in_buf[448]*(-6)+in_buf[449]*(-16)+in_buf[450]*(-2)+in_buf[451]*(-4)+in_buf[452]*(-7)+in_buf[453]*(-15)+in_buf[454]*(-8)+in_buf[455]*(0)+in_buf[456]*(15)+in_buf[457]*(-3)+in_buf[458]*(2)+in_buf[459]*(2)+in_buf[460]*(1)+in_buf[461]*(-1)+in_buf[462]*(-5)+in_buf[463]*(-6)+in_buf[464]*(-11)+in_buf[465]*(-1)+in_buf[466]*(-13)+in_buf[467]*(-23)+in_buf[468]*(1)+in_buf[469]*(-6)+in_buf[470]*(5)+in_buf[471]*(14)+in_buf[472]*(3)+in_buf[473]*(16)+in_buf[474]*(-35)+in_buf[475]*(-30)+in_buf[476]*(1)+in_buf[477]*(-8)+in_buf[478]*(-8)+in_buf[479]*(-4)+in_buf[480]*(4)+in_buf[481]*(0)+in_buf[482]*(4)+in_buf[483]*(-4)+in_buf[484]*(3)+in_buf[485]*(8)+in_buf[486]*(0)+in_buf[487]*(-2)+in_buf[488]*(-7)+in_buf[489]*(-7)+in_buf[490]*(-14)+in_buf[491]*(-10)+in_buf[492]*(-7)+in_buf[493]*(7)+in_buf[494]*(-14)+in_buf[495]*(-11)+in_buf[496]*(11)+in_buf[497]*(5)+in_buf[498]*(12)+in_buf[499]*(22)+in_buf[500]*(24)+in_buf[501]*(-14)+in_buf[502]*(-25)+in_buf[503]*(7)+in_buf[504]*(-30)+in_buf[505]*(-15)+in_buf[506]*(-24)+in_buf[507]*(-17)+in_buf[508]*(1)+in_buf[509]*(11)+in_buf[510]*(14)+in_buf[511]*(5)+in_buf[512]*(5)+in_buf[513]*(1)+in_buf[514]*(0)+in_buf[515]*(-3)+in_buf[516]*(-1)+in_buf[517]*(-18)+in_buf[518]*(-11)+in_buf[519]*(-2)+in_buf[520]*(-4)+in_buf[521]*(-11)+in_buf[522]*(-16)+in_buf[523]*(-12)+in_buf[524]*(6)+in_buf[525]*(7)+in_buf[526]*(8)+in_buf[527]*(6)+in_buf[528]*(1)+in_buf[529]*(-24)+in_buf[530]*(-31)+in_buf[531]*(-23)+in_buf[532]*(-20)+in_buf[533]*(-4)+in_buf[534]*(-10)+in_buf[535]*(-14)+in_buf[536]*(-1)+in_buf[537]*(11)+in_buf[538]*(13)+in_buf[539]*(1)+in_buf[540]*(14)+in_buf[541]*(1)+in_buf[542]*(4)+in_buf[543]*(-5)+in_buf[544]*(1)+in_buf[545]*(-7)+in_buf[546]*(-4)+in_buf[547]*(0)+in_buf[548]*(-4)+in_buf[549]*(-5)+in_buf[550]*(-5)+in_buf[551]*(-6)+in_buf[552]*(15)+in_buf[553]*(8)+in_buf[554]*(10)+in_buf[555]*(3)+in_buf[556]*(0)+in_buf[557]*(-38)+in_buf[558]*(-23)+in_buf[559]*(-11)+in_buf[560]*(-1)+in_buf[561]*(28)+in_buf[562]*(-4)+in_buf[563]*(-24)+in_buf[564]*(3)+in_buf[565]*(14)+in_buf[566]*(-1)+in_buf[567]*(1)+in_buf[568]*(22)+in_buf[569]*(14)+in_buf[570]*(14)+in_buf[571]*(7)+in_buf[572]*(10)+in_buf[573]*(12)+in_buf[574]*(-2)+in_buf[575]*(1)+in_buf[576]*(-8)+in_buf[577]*(-6)+in_buf[578]*(-17)+in_buf[579]*(1)+in_buf[580]*(15)+in_buf[581]*(12)+in_buf[582]*(10)+in_buf[583]*(-7)+in_buf[584]*(-15)+in_buf[585]*(-3)+in_buf[586]*(-25)+in_buf[587]*(-6)+in_buf[588]*(-22)+in_buf[589]*(-6)+in_buf[590]*(-27)+in_buf[591]*(-15)+in_buf[592]*(11)+in_buf[593]*(8)+in_buf[594]*(5)+in_buf[595]*(6)+in_buf[596]*(10)+in_buf[597]*(13)+in_buf[598]*(4)+in_buf[599]*(21)+in_buf[600]*(9)+in_buf[601]*(10)+in_buf[602]*(4)+in_buf[603]*(16)+in_buf[604]*(-1)+in_buf[605]*(3)+in_buf[606]*(-14)+in_buf[607]*(-10)+in_buf[608]*(-4)+in_buf[609]*(-3)+in_buf[610]*(3)+in_buf[611]*(-12)+in_buf[612]*(-25)+in_buf[613]*(-8)+in_buf[614]*(32)+in_buf[615]*(2)+in_buf[616]*(-23)+in_buf[617]*(-13)+in_buf[618]*(-43)+in_buf[619]*(-6)+in_buf[620]*(1)+in_buf[621]*(-14)+in_buf[622]*(13)+in_buf[623]*(17)+in_buf[624]*(4)+in_buf[625]*(7)+in_buf[626]*(5)+in_buf[627]*(21)+in_buf[628]*(26)+in_buf[629]*(16)+in_buf[630]*(18)+in_buf[631]*(14)+in_buf[632]*(12)+in_buf[633]*(5)+in_buf[634]*(-18)+in_buf[635]*(-15)+in_buf[636]*(-23)+in_buf[637]*(-15)+in_buf[638]*(1)+in_buf[639]*(3)+in_buf[640]*(-26)+in_buf[641]*(0)+in_buf[642]*(22)+in_buf[643]*(4)+in_buf[644]*(1)+in_buf[645]*(4)+in_buf[646]*(-32)+in_buf[647]*(23)+in_buf[648]*(12)+in_buf[649]*(-7)+in_buf[650]*(-10)+in_buf[651]*(-1)+in_buf[652]*(22)+in_buf[653]*(6)+in_buf[654]*(11)+in_buf[655]*(9)+in_buf[656]*(6)+in_buf[657]*(8)+in_buf[658]*(17)+in_buf[659]*(19)+in_buf[660]*(17)+in_buf[661]*(2)+in_buf[662]*(1)+in_buf[663]*(-15)+in_buf[664]*(-16)+in_buf[665]*(-2)+in_buf[666]*(-6)+in_buf[667]*(-3)+in_buf[668]*(-23)+in_buf[669]*(1)+in_buf[670]*(-8)+in_buf[671]*(3)+in_buf[672]*(-1)+in_buf[673]*(0)+in_buf[674]*(-16)+in_buf[675]*(1)+in_buf[676]*(-30)+in_buf[677]*(4)+in_buf[678]*(-2)+in_buf[679]*(-2)+in_buf[680]*(-1)+in_buf[681]*(6)+in_buf[682]*(4)+in_buf[683]*(1)+in_buf[684]*(20)+in_buf[685]*(23)+in_buf[686]*(15)+in_buf[687]*(20)+in_buf[688]*(8)+in_buf[689]*(-31)+in_buf[690]*(-7)+in_buf[691]*(0)+in_buf[692]*(1)+in_buf[693]*(-38)+in_buf[694]*(-16)+in_buf[695]*(-8)+in_buf[696]*(-22)+in_buf[697]*(-22)+in_buf[698]*(-19)+in_buf[699]*(4)+in_buf[700]*(0)+in_buf[701]*(-1)+in_buf[702]*(25)+in_buf[703]*(0)+in_buf[704]*(-25)+in_buf[705]*(-17)+in_buf[706]*(-12)+in_buf[707]*(-11)+in_buf[708]*(-37)+in_buf[709]*(-18)+in_buf[710]*(12)+in_buf[711]*(-1)+in_buf[712]*(-19)+in_buf[713]*(0)+in_buf[714]*(-18)+in_buf[715]*(1)+in_buf[716]*(-9)+in_buf[717]*(-7)+in_buf[718]*(-2)+in_buf[719]*(30)+in_buf[720]*(17)+in_buf[721]*(8)+in_buf[722]*(9)+in_buf[723]*(16)+in_buf[724]*(21)+in_buf[725]*(-2)+in_buf[726]*(-10)+in_buf[727]*(2)+in_buf[728]*(-2)+in_buf[729]*(0)+in_buf[730]*(-2)+in_buf[731]*(17)+in_buf[732]*(42)+in_buf[733]*(39)+in_buf[734]*(16)+in_buf[735]*(-17)+in_buf[736]*(6)+in_buf[737]*(-12)+in_buf[738]*(-8)+in_buf[739]*(4)+in_buf[740]*(23)+in_buf[741]*(4)+in_buf[742]*(0)+in_buf[743]*(-10)+in_buf[744]*(-2)+in_buf[745]*(-3)+in_buf[746]*(1)+in_buf[747]*(-6)+in_buf[748]*(-3)+in_buf[749]*(-15)+in_buf[750]*(-5)+in_buf[751]*(17)+in_buf[752]*(8)+in_buf[753]*(-12)+in_buf[754]*(-3)+in_buf[755]*(2)+in_buf[756]*(1)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(-1)+in_buf[760]*(-22)+in_buf[761]*(-17)+in_buf[762]*(3)+in_buf[763]*(4)+in_buf[764]*(4)+in_buf[765]*(-11)+in_buf[766]*(11)+in_buf[767]*(0)+in_buf[768]*(1)+in_buf[769]*(-20)+in_buf[770]*(-9)+in_buf[771]*(0)+in_buf[772]*(-17)+in_buf[773]*(-32)+in_buf[774]*(-23)+in_buf[775]*(11)+in_buf[776]*(12)+in_buf[777]*(-21)+in_buf[778]*(-27)+in_buf[779]*(-23)+in_buf[780]*(-2)+in_buf[781]*(0)+in_buf[782]*(-1)+in_buf[783]*(-2);
assign in_buf_weight040=in_buf[0]*(-3)+in_buf[1]*(0)+in_buf[2]*(3)+in_buf[3]*(4)+in_buf[4]*(-1)+in_buf[5]*(2)+in_buf[6]*(0)+in_buf[7]*(1)+in_buf[8]*(4)+in_buf[9]*(1)+in_buf[10]*(-2)+in_buf[11]*(0)+in_buf[12]*(-9)+in_buf[13]*(-5)+in_buf[14]*(14)+in_buf[15]*(12)+in_buf[16]*(4)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(-2)+in_buf[20]*(2)+in_buf[21]*(-3)+in_buf[22]*(3)+in_buf[23]*(-1)+in_buf[24]*(1)+in_buf[25]*(0)+in_buf[26]*(0)+in_buf[27]*(-2)+in_buf[28]*(2)+in_buf[29]*(4)+in_buf[30]*(0)+in_buf[31]*(-1)+in_buf[32]*(2)+in_buf[33]*(4)+in_buf[34]*(14)+in_buf[35]*(2)+in_buf[36]*(2)+in_buf[37]*(-3)+in_buf[38]*(-17)+in_buf[39]*(-11)+in_buf[40]*(-2)+in_buf[41]*(-4)+in_buf[42]*(0)+in_buf[43]*(10)+in_buf[44]*(21)+in_buf[45]*(-3)+in_buf[46]*(-15)+in_buf[47]*(-14)+in_buf[48]*(-3)+in_buf[49]*(-6)+in_buf[50]*(0)+in_buf[51]*(1)+in_buf[52]*(0)+in_buf[53]*(0)+in_buf[54]*(3)+in_buf[55]*(3)+in_buf[56]*(1)+in_buf[57]*(-1)+in_buf[58]*(-1)+in_buf[59]*(10)+in_buf[60]*(-1)+in_buf[61]*(-4)+in_buf[62]*(-7)+in_buf[63]*(-3)+in_buf[64]*(4)+in_buf[65]*(29)+in_buf[66]*(28)+in_buf[67]*(20)+in_buf[68]*(-11)+in_buf[69]*(-8)+in_buf[70]*(-6)+in_buf[71]*(-35)+in_buf[72]*(-39)+in_buf[73]*(-31)+in_buf[74]*(-38)+in_buf[75]*(-38)+in_buf[76]*(-31)+in_buf[77]*(-9)+in_buf[78]*(-7)+in_buf[79]*(2)+in_buf[80]*(1)+in_buf[81]*(4)+in_buf[82]*(0)+in_buf[83]*(-1)+in_buf[84]*(-1)+in_buf[85]*(1)+in_buf[86]*(21)+in_buf[87]*(6)+in_buf[88]*(-3)+in_buf[89]*(-2)+in_buf[90]*(12)+in_buf[91]*(33)+in_buf[92]*(58)+in_buf[93]*(46)+in_buf[94]*(44)+in_buf[95]*(29)+in_buf[96]*(8)+in_buf[97]*(4)+in_buf[98]*(0)+in_buf[99]*(-38)+in_buf[100]*(-32)+in_buf[101]*(-14)+in_buf[102]*(-23)+in_buf[103]*(-29)+in_buf[104]*(-16)+in_buf[105]*(-16)+in_buf[106]*(-30)+in_buf[107]*(-25)+in_buf[108]*(-9)+in_buf[109]*(0)+in_buf[110]*(-7)+in_buf[111]*(-3)+in_buf[112]*(0)+in_buf[113]*(4)+in_buf[114]*(26)+in_buf[115]*(35)+in_buf[116]*(46)+in_buf[117]*(14)+in_buf[118]*(6)+in_buf[119]*(0)+in_buf[120]*(23)+in_buf[121]*(19)+in_buf[122]*(6)+in_buf[123]*(20)+in_buf[124]*(16)+in_buf[125]*(-4)+in_buf[126]*(-3)+in_buf[127]*(-14)+in_buf[128]*(-23)+in_buf[129]*(-8)+in_buf[130]*(3)+in_buf[131]*(-5)+in_buf[132]*(-24)+in_buf[133]*(-51)+in_buf[134]*(-52)+in_buf[135]*(-37)+in_buf[136]*(-25)+in_buf[137]*(-9)+in_buf[138]*(-2)+in_buf[139]*(0)+in_buf[140]*(0)+in_buf[141]*(4)+in_buf[142]*(-5)+in_buf[143]*(18)+in_buf[144]*(37)+in_buf[145]*(32)+in_buf[146]*(14)+in_buf[147]*(1)+in_buf[148]*(7)+in_buf[149]*(12)+in_buf[150]*(12)+in_buf[151]*(25)+in_buf[152]*(27)+in_buf[153]*(29)+in_buf[154]*(28)+in_buf[155]*(27)+in_buf[156]*(14)+in_buf[157]*(9)+in_buf[158]*(-6)+in_buf[159]*(-14)+in_buf[160]*(-30)+in_buf[161]*(-36)+in_buf[162]*(-54)+in_buf[163]*(-37)+in_buf[164]*(-21)+in_buf[165]*(-7)+in_buf[166]*(0)+in_buf[167]*(-3)+in_buf[168]*(-3)+in_buf[169]*(23)+in_buf[170]*(27)+in_buf[171]*(59)+in_buf[172]*(36)+in_buf[173]*(22)+in_buf[174]*(23)+in_buf[175]*(2)+in_buf[176]*(2)+in_buf[177]*(21)+in_buf[178]*(48)+in_buf[179]*(37)+in_buf[180]*(41)+in_buf[181]*(48)+in_buf[182]*(55)+in_buf[183]*(61)+in_buf[184]*(40)+in_buf[185]*(20)+in_buf[186]*(3)+in_buf[187]*(-6)+in_buf[188]*(-10)+in_buf[189]*(-14)+in_buf[190]*(-26)+in_buf[191]*(-33)+in_buf[192]*(-54)+in_buf[193]*(-29)+in_buf[194]*(5)+in_buf[195]*(-10)+in_buf[196]*(0)+in_buf[197]*(33)+in_buf[198]*(39)+in_buf[199]*(74)+in_buf[200]*(12)+in_buf[201]*(-1)+in_buf[202]*(13)+in_buf[203]*(4)+in_buf[204]*(18)+in_buf[205]*(23)+in_buf[206]*(32)+in_buf[207]*(41)+in_buf[208]*(44)+in_buf[209]*(53)+in_buf[210]*(65)+in_buf[211]*(48)+in_buf[212]*(19)+in_buf[213]*(6)+in_buf[214]*(0)+in_buf[215]*(-11)+in_buf[216]*(-13)+in_buf[217]*(-22)+in_buf[218]*(-27)+in_buf[219]*(-55)+in_buf[220]*(-61)+in_buf[221]*(-39)+in_buf[222]*(-11)+in_buf[223]*(-4)+in_buf[224]*(12)+in_buf[225]*(31)+in_buf[226]*(41)+in_buf[227]*(36)+in_buf[228]*(5)+in_buf[229]*(11)+in_buf[230]*(7)+in_buf[231]*(15)+in_buf[232]*(31)+in_buf[233]*(25)+in_buf[234]*(32)+in_buf[235]*(21)+in_buf[236]*(24)+in_buf[237]*(22)+in_buf[238]*(33)+in_buf[239]*(12)+in_buf[240]*(-3)+in_buf[241]*(-11)+in_buf[242]*(13)+in_buf[243]*(5)+in_buf[244]*(-2)+in_buf[245]*(-10)+in_buf[246]*(-9)+in_buf[247]*(-54)+in_buf[248]*(-70)+in_buf[249]*(-41)+in_buf[250]*(-20)+in_buf[251]*(7)+in_buf[252]*(6)+in_buf[253]*(16)+in_buf[254]*(51)+in_buf[255]*(19)+in_buf[256]*(7)+in_buf[257]*(4)+in_buf[258]*(19)+in_buf[259]*(16)+in_buf[260]*(29)+in_buf[261]*(34)+in_buf[262]*(13)+in_buf[263]*(-9)+in_buf[264]*(-4)+in_buf[265]*(-20)+in_buf[266]*(-23)+in_buf[267]*(-24)+in_buf[268]*(-19)+in_buf[269]*(11)+in_buf[270]*(18)+in_buf[271]*(23)+in_buf[272]*(9)+in_buf[273]*(0)+in_buf[274]*(-4)+in_buf[275]*(-41)+in_buf[276]*(-63)+in_buf[277]*(-32)+in_buf[278]*(-1)+in_buf[279]*(6)+in_buf[280]*(13)+in_buf[281]*(11)+in_buf[282]*(39)+in_buf[283]*(22)+in_buf[284]*(-18)+in_buf[285]*(-6)+in_buf[286]*(23)+in_buf[287]*(22)+in_buf[288]*(14)+in_buf[289]*(2)+in_buf[290]*(-19)+in_buf[291]*(-35)+in_buf[292]*(-63)+in_buf[293]*(-58)+in_buf[294]*(-37)+in_buf[295]*(-32)+in_buf[296]*(0)+in_buf[297]*(17)+in_buf[298]*(32)+in_buf[299]*(13)+in_buf[300]*(14)+in_buf[301]*(25)+in_buf[302]*(15)+in_buf[303]*(-13)+in_buf[304]*(-48)+in_buf[305]*(-44)+in_buf[306]*(-18)+in_buf[307]*(9)+in_buf[308]*(17)+in_buf[309]*(2)+in_buf[310]*(20)+in_buf[311]*(-6)+in_buf[312]*(-17)+in_buf[313]*(0)+in_buf[314]*(17)+in_buf[315]*(-1)+in_buf[316]*(-9)+in_buf[317]*(-10)+in_buf[318]*(-24)+in_buf[319]*(-36)+in_buf[320]*(-44)+in_buf[321]*(-33)+in_buf[322]*(-16)+in_buf[323]*(-5)+in_buf[324]*(3)+in_buf[325]*(31)+in_buf[326]*(18)+in_buf[327]*(13)+in_buf[328]*(22)+in_buf[329]*(20)+in_buf[330]*(21)+in_buf[331]*(6)+in_buf[332]*(-23)+in_buf[333]*(-44)+in_buf[334]*(-20)+in_buf[335]*(-24)+in_buf[336]*(16)+in_buf[337]*(-2)+in_buf[338]*(8)+in_buf[339]*(12)+in_buf[340]*(5)+in_buf[341]*(-3)+in_buf[342]*(0)+in_buf[343]*(-30)+in_buf[344]*(-25)+in_buf[345]*(-25)+in_buf[346]*(-33)+in_buf[347]*(-39)+in_buf[348]*(-39)+in_buf[349]*(-10)+in_buf[350]*(9)+in_buf[351]*(10)+in_buf[352]*(7)+in_buf[353]*(8)+in_buf[354]*(6)+in_buf[355]*(7)+in_buf[356]*(7)+in_buf[357]*(15)+in_buf[358]*(2)+in_buf[359]*(15)+in_buf[360]*(-29)+in_buf[361]*(-31)+in_buf[362]*(-5)+in_buf[363]*(-4)+in_buf[364]*(-18)+in_buf[365]*(-4)+in_buf[366]*(-3)+in_buf[367]*(24)+in_buf[368]*(-6)+in_buf[369]*(-30)+in_buf[370]*(-23)+in_buf[371]*(-20)+in_buf[372]*(-15)+in_buf[373]*(-10)+in_buf[374]*(-3)+in_buf[375]*(-24)+in_buf[376]*(-16)+in_buf[377]*(-6)+in_buf[378]*(-9)+in_buf[379]*(-1)+in_buf[380]*(11)+in_buf[381]*(-1)+in_buf[382]*(-3)+in_buf[383]*(-9)+in_buf[384]*(2)+in_buf[385]*(12)+in_buf[386]*(6)+in_buf[387]*(2)+in_buf[388]*(-23)+in_buf[389]*(-38)+in_buf[390]*(-4)+in_buf[391]*(12)+in_buf[392]*(-18)+in_buf[393]*(4)+in_buf[394]*(-6)+in_buf[395]*(5)+in_buf[396]*(-6)+in_buf[397]*(-37)+in_buf[398]*(-23)+in_buf[399]*(-6)+in_buf[400]*(-6)+in_buf[401]*(-9)+in_buf[402]*(-4)+in_buf[403]*(-15)+in_buf[404]*(-6)+in_buf[405]*(0)+in_buf[406]*(-11)+in_buf[407]*(3)+in_buf[408]*(-1)+in_buf[409]*(-1)+in_buf[410]*(7)+in_buf[411]*(-5)+in_buf[412]*(2)+in_buf[413]*(14)+in_buf[414]*(11)+in_buf[415]*(-1)+in_buf[416]*(-9)+in_buf[417]*(-15)+in_buf[418]*(2)+in_buf[419]*(10)+in_buf[420]*(-18)+in_buf[421]*(15)+in_buf[422]*(-11)+in_buf[423]*(-21)+in_buf[424]*(2)+in_buf[425]*(-15)+in_buf[426]*(-5)+in_buf[427]*(-9)+in_buf[428]*(-10)+in_buf[429]*(-17)+in_buf[430]*(-17)+in_buf[431]*(-16)+in_buf[432]*(-15)+in_buf[433]*(-16)+in_buf[434]*(-5)+in_buf[435]*(10)+in_buf[436]*(-7)+in_buf[437]*(0)+in_buf[438]*(-5)+in_buf[439]*(-20)+in_buf[440]*(-3)+in_buf[441]*(12)+in_buf[442]*(15)+in_buf[443]*(-9)+in_buf[444]*(0)+in_buf[445]*(-4)+in_buf[446]*(-9)+in_buf[447]*(29)+in_buf[448]*(0)+in_buf[449]*(29)+in_buf[450]*(15)+in_buf[451]*(-7)+in_buf[452]*(14)+in_buf[453]*(0)+in_buf[454]*(-10)+in_buf[455]*(-17)+in_buf[456]*(-24)+in_buf[457]*(-20)+in_buf[458]*(-15)+in_buf[459]*(-9)+in_buf[460]*(-1)+in_buf[461]*(2)+in_buf[462]*(4)+in_buf[463]*(-8)+in_buf[464]*(-7)+in_buf[465]*(0)+in_buf[466]*(-8)+in_buf[467]*(-16)+in_buf[468]*(0)+in_buf[469]*(-3)+in_buf[470]*(11)+in_buf[471]*(-2)+in_buf[472]*(-2)+in_buf[473]*(-12)+in_buf[474]*(-8)+in_buf[475]*(23)+in_buf[476]*(-2)+in_buf[477]*(14)+in_buf[478]*(-5)+in_buf[479]*(28)+in_buf[480]*(35)+in_buf[481]*(4)+in_buf[482]*(-21)+in_buf[483]*(-27)+in_buf[484]*(-35)+in_buf[485]*(-21)+in_buf[486]*(-5)+in_buf[487]*(-2)+in_buf[488]*(9)+in_buf[489]*(6)+in_buf[490]*(-7)+in_buf[491]*(-1)+in_buf[492]*(-3)+in_buf[493]*(7)+in_buf[494]*(-11)+in_buf[495]*(-1)+in_buf[496]*(2)+in_buf[497]*(-20)+in_buf[498]*(-6)+in_buf[499]*(-19)+in_buf[500]*(-13)+in_buf[501]*(28)+in_buf[502]*(8)+in_buf[503]*(-2)+in_buf[504]*(13)+in_buf[505]*(6)+in_buf[506]*(-7)+in_buf[507]*(26)+in_buf[508]*(18)+in_buf[509]*(17)+in_buf[510]*(-4)+in_buf[511]*(-23)+in_buf[512]*(-33)+in_buf[513]*(-15)+in_buf[514]*(18)+in_buf[515]*(16)+in_buf[516]*(12)+in_buf[517]*(0)+in_buf[518]*(-13)+in_buf[519]*(-4)+in_buf[520]*(3)+in_buf[521]*(14)+in_buf[522]*(7)+in_buf[523]*(27)+in_buf[524]*(8)+in_buf[525]*(-6)+in_buf[526]*(1)+in_buf[527]*(-12)+in_buf[528]*(-5)+in_buf[529]*(28)+in_buf[530]*(38)+in_buf[531]*(3)+in_buf[532]*(-20)+in_buf[533]*(7)+in_buf[534]*(-9)+in_buf[535]*(11)+in_buf[536]*(16)+in_buf[537]*(10)+in_buf[538]*(-17)+in_buf[539]*(-15)+in_buf[540]*(-16)+in_buf[541]*(-1)+in_buf[542]*(28)+in_buf[543]*(19)+in_buf[544]*(20)+in_buf[545]*(-5)+in_buf[546]*(-14)+in_buf[547]*(-1)+in_buf[548]*(15)+in_buf[549]*(6)+in_buf[550]*(13)+in_buf[551]*(26)+in_buf[552]*(11)+in_buf[553]*(-7)+in_buf[554]*(-1)+in_buf[555]*(-19)+in_buf[556]*(5)+in_buf[557]*(4)+in_buf[558]*(8)+in_buf[559]*(8)+in_buf[560]*(0)+in_buf[561]*(24)+in_buf[562]*(-19)+in_buf[563]*(-6)+in_buf[564]*(13)+in_buf[565]*(19)+in_buf[566]*(-17)+in_buf[567]*(-14)+in_buf[568]*(-15)+in_buf[569]*(-2)+in_buf[570]*(8)+in_buf[571]*(2)+in_buf[572]*(-9)+in_buf[573]*(-5)+in_buf[574]*(-3)+in_buf[575]*(0)+in_buf[576]*(13)+in_buf[577]*(1)+in_buf[578]*(1)+in_buf[579]*(22)+in_buf[580]*(9)+in_buf[581]*(-7)+in_buf[582]*(-16)+in_buf[583]*(-10)+in_buf[584]*(30)+in_buf[585]*(10)+in_buf[586]*(-11)+in_buf[587]*(-9)+in_buf[588]*(-17)+in_buf[589]*(11)+in_buf[590]*(21)+in_buf[591]*(-29)+in_buf[592]*(2)+in_buf[593]*(-9)+in_buf[594]*(-25)+in_buf[595]*(-16)+in_buf[596]*(-28)+in_buf[597]*(-29)+in_buf[598]*(-11)+in_buf[599]*(-11)+in_buf[600]*(2)+in_buf[601]*(0)+in_buf[602]*(5)+in_buf[603]*(0)+in_buf[604]*(20)+in_buf[605]*(2)+in_buf[606]*(1)+in_buf[607]*(9)+in_buf[608]*(14)+in_buf[609]*(-3)+in_buf[610]*(-20)+in_buf[611]*(-18)+in_buf[612]*(16)+in_buf[613]*(-21)+in_buf[614]*(18)+in_buf[615]*(6)+in_buf[616]*(-15)+in_buf[617]*(12)+in_buf[618]*(27)+in_buf[619]*(-26)+in_buf[620]*(1)+in_buf[621]*(0)+in_buf[622]*(-2)+in_buf[623]*(-7)+in_buf[624]*(-20)+in_buf[625]*(-23)+in_buf[626]*(-13)+in_buf[627]*(-2)+in_buf[628]*(13)+in_buf[629]*(10)+in_buf[630]*(22)+in_buf[631]*(7)+in_buf[632]*(25)+in_buf[633]*(5)+in_buf[634]*(-9)+in_buf[635]*(-11)+in_buf[636]*(2)+in_buf[637]*(-19)+in_buf[638]*(-14)+in_buf[639]*(-9)+in_buf[640]*(28)+in_buf[641]*(-31)+in_buf[642]*(-11)+in_buf[643]*(4)+in_buf[644]*(0)+in_buf[645]*(3)+in_buf[646]*(40)+in_buf[647]*(-22)+in_buf[648]*(-20)+in_buf[649]*(6)+in_buf[650]*(9)+in_buf[651]*(7)+in_buf[652]*(-10)+in_buf[653]*(-3)+in_buf[654]*(0)+in_buf[655]*(38)+in_buf[656]*(14)+in_buf[657]*(0)+in_buf[658]*(14)+in_buf[659]*(22)+in_buf[660]*(9)+in_buf[661]*(7)+in_buf[662]*(5)+in_buf[663]*(-5)+in_buf[664]*(10)+in_buf[665]*(-9)+in_buf[666]*(9)+in_buf[667]*(9)+in_buf[668]*(23)+in_buf[669]*(-19)+in_buf[670]*(-34)+in_buf[671]*(-2)+in_buf[672]*(2)+in_buf[673]*(2)+in_buf[674]*(24)+in_buf[675]*(28)+in_buf[676]*(58)+in_buf[677]*(47)+in_buf[678]*(20)+in_buf[679]*(20)+in_buf[680]*(14)+in_buf[681]*(14)+in_buf[682]*(25)+in_buf[683]*(17)+in_buf[684]*(7)+in_buf[685]*(10)+in_buf[686]*(10)+in_buf[687]*(20)+in_buf[688]*(12)+in_buf[689]*(8)+in_buf[690]*(-4)+in_buf[691]*(-13)+in_buf[692]*(3)+in_buf[693]*(-9)+in_buf[694]*(4)+in_buf[695]*(27)+in_buf[696]*(1)+in_buf[697]*(-20)+in_buf[698]*(-14)+in_buf[699]*(1)+in_buf[700]*(-3)+in_buf[701]*(0)+in_buf[702]*(22)+in_buf[703]*(5)+in_buf[704]*(4)+in_buf[705]*(7)+in_buf[706]*(-5)+in_buf[707]*(5)+in_buf[708]*(36)+in_buf[709]*(39)+in_buf[710]*(56)+in_buf[711]*(33)+in_buf[712]*(13)+in_buf[713]*(12)+in_buf[714]*(14)+in_buf[715]*(6)+in_buf[716]*(5)+in_buf[717]*(-15)+in_buf[718]*(1)+in_buf[719]*(13)+in_buf[720]*(7)+in_buf[721]*(16)+in_buf[722]*(2)+in_buf[723]*(11)+in_buf[724]*(14)+in_buf[725]*(-7)+in_buf[726]*(-3)+in_buf[727]*(2)+in_buf[728]*(0)+in_buf[729]*(3)+in_buf[730]*(3)+in_buf[731]*(8)+in_buf[732]*(-18)+in_buf[733]*(-24)+in_buf[734]*(-13)+in_buf[735]*(24)+in_buf[736]*(27)+in_buf[737]*(30)+in_buf[738]*(29)+in_buf[739]*(36)+in_buf[740]*(29)+in_buf[741]*(45)+in_buf[742]*(34)+in_buf[743]*(1)+in_buf[744]*(24)+in_buf[745]*(40)+in_buf[746]*(66)+in_buf[747]*(46)+in_buf[748]*(50)+in_buf[749]*(21)+in_buf[750]*(40)+in_buf[751]*(20)+in_buf[752]*(-11)+in_buf[753]*(11)+in_buf[754]*(4)+in_buf[755]*(4)+in_buf[756]*(2)+in_buf[757]*(-2)+in_buf[758]*(2)+in_buf[759]*(2)+in_buf[760]*(6)+in_buf[761]*(16)+in_buf[762]*(11)+in_buf[763]*(9)+in_buf[764]*(11)+in_buf[765]*(3)+in_buf[766]*(37)+in_buf[767]*(9)+in_buf[768]*(1)+in_buf[769]*(-14)+in_buf[770]*(0)+in_buf[771]*(-4)+in_buf[772]*(4)+in_buf[773]*(-1)+in_buf[774]*(7)+in_buf[775]*(41)+in_buf[776]*(40)+in_buf[777]*(34)+in_buf[778]*(16)+in_buf[779]*(5)+in_buf[780]*(3)+in_buf[781]*(-2)+in_buf[782]*(-2)+in_buf[783]*(0);
assign in_buf_weight041=in_buf[0]*(2)+in_buf[1]*(0)+in_buf[2]*(4)+in_buf[3]*(3)+in_buf[4]*(0)+in_buf[5]*(0)+in_buf[6]*(0)+in_buf[7]*(0)+in_buf[8]*(-1)+in_buf[9]*(3)+in_buf[10]*(0)+in_buf[11]*(4)+in_buf[12]*(11)+in_buf[13]*(12)+in_buf[14]*(-9)+in_buf[15]*(-4)+in_buf[16]*(4)+in_buf[17]*(2)+in_buf[18]*(-1)+in_buf[19]*(0)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(-3)+in_buf[23]*(1)+in_buf[24]*(2)+in_buf[25]*(0)+in_buf[26]*(-2)+in_buf[27]*(-1)+in_buf[28]*(2)+in_buf[29]*(1)+in_buf[30]*(-1)+in_buf[31]*(-2)+in_buf[32]*(4)+in_buf[33]*(-4)+in_buf[34]*(-4)+in_buf[35]*(-4)+in_buf[36]*(9)+in_buf[37]*(11)+in_buf[38]*(32)+in_buf[39]*(8)+in_buf[40]*(-7)+in_buf[41]*(10)+in_buf[42]*(11)+in_buf[43]*(-8)+in_buf[44]*(-23)+in_buf[45]*(-4)+in_buf[46]*(19)+in_buf[47]*(27)+in_buf[48]*(36)+in_buf[49]*(25)+in_buf[50]*(20)+in_buf[51]*(13)+in_buf[52]*(2)+in_buf[53]*(-1)+in_buf[54]*(3)+in_buf[55]*(0)+in_buf[56]*(-3)+in_buf[57]*(2)+in_buf[58]*(12)+in_buf[59]*(-28)+in_buf[60]*(-21)+in_buf[61]*(7)+in_buf[62]*(5)+in_buf[63]*(14)+in_buf[64]*(9)+in_buf[65]*(0)+in_buf[66]*(-9)+in_buf[67]*(-13)+in_buf[68]*(-2)+in_buf[69]*(31)+in_buf[70]*(31)+in_buf[71]*(18)+in_buf[72]*(-7)+in_buf[73]*(14)+in_buf[74]*(23)+in_buf[75]*(17)+in_buf[76]*(8)+in_buf[77]*(17)+in_buf[78]*(61)+in_buf[79]*(25)+in_buf[80]*(-2)+in_buf[81]*(-2)+in_buf[82]*(-2)+in_buf[83]*(1)+in_buf[84]*(-1)+in_buf[85]*(4)+in_buf[86]*(-2)+in_buf[87]*(-31)+in_buf[88]*(-14)+in_buf[89]*(-7)+in_buf[90]*(17)+in_buf[91]*(21)+in_buf[92]*(5)+in_buf[93]*(15)+in_buf[94]*(14)+in_buf[95]*(11)+in_buf[96]*(1)+in_buf[97]*(1)+in_buf[98]*(-18)+in_buf[99]*(-21)+in_buf[100]*(-21)+in_buf[101]*(-14)+in_buf[102]*(-11)+in_buf[103]*(-8)+in_buf[104]*(-4)+in_buf[105]*(22)+in_buf[106]*(54)+in_buf[107]*(65)+in_buf[108]*(10)+in_buf[109]*(-23)+in_buf[110]*(-3)+in_buf[111]*(-3)+in_buf[112]*(0)+in_buf[113]*(1)+in_buf[114]*(-10)+in_buf[115]*(-1)+in_buf[116]*(5)+in_buf[117]*(-6)+in_buf[118]*(-2)+in_buf[119]*(21)+in_buf[120]*(3)+in_buf[121]*(10)+in_buf[122]*(13)+in_buf[123]*(4)+in_buf[124]*(-6)+in_buf[125]*(-1)+in_buf[126]*(11)+in_buf[127]*(4)+in_buf[128]*(1)+in_buf[129]*(7)+in_buf[130]*(-1)+in_buf[131]*(7)+in_buf[132]*(19)+in_buf[133]*(35)+in_buf[134]*(34)+in_buf[135]*(66)+in_buf[136]*(59)+in_buf[137]*(28)+in_buf[138]*(-34)+in_buf[139]*(2)+in_buf[140]*(0)+in_buf[141]*(-1)+in_buf[142]*(11)+in_buf[143]*(-29)+in_buf[144]*(-46)+in_buf[145]*(-8)+in_buf[146]*(1)+in_buf[147]*(13)+in_buf[148]*(5)+in_buf[149]*(14)+in_buf[150]*(17)+in_buf[151]*(-7)+in_buf[152]*(-9)+in_buf[153]*(-13)+in_buf[154]*(1)+in_buf[155]*(-9)+in_buf[156]*(-16)+in_buf[157]*(-20)+in_buf[158]*(-13)+in_buf[159]*(-2)+in_buf[160]*(17)+in_buf[161]*(23)+in_buf[162]*(2)+in_buf[163]*(19)+in_buf[164]*(42)+in_buf[165]*(23)+in_buf[166]*(-14)+in_buf[167]*(11)+in_buf[168]*(3)+in_buf[169]*(-5)+in_buf[170]*(-7)+in_buf[171]*(-35)+in_buf[172]*(-16)+in_buf[173]*(14)+in_buf[174]*(0)+in_buf[175]*(14)+in_buf[176]*(17)+in_buf[177]*(18)+in_buf[178]*(-12)+in_buf[179]*(-5)+in_buf[180]*(-7)+in_buf[181]*(-18)+in_buf[182]*(-8)+in_buf[183]*(-7)+in_buf[184]*(-25)+in_buf[185]*(-1)+in_buf[186]*(-11)+in_buf[187]*(5)+in_buf[188]*(18)+in_buf[189]*(-3)+in_buf[190]*(-13)+in_buf[191]*(0)+in_buf[192]*(13)+in_buf[193]*(21)+in_buf[194]*(15)+in_buf[195]*(14)+in_buf[196]*(5)+in_buf[197]*(-11)+in_buf[198]*(-4)+in_buf[199]*(-17)+in_buf[200]*(-26)+in_buf[201]*(3)+in_buf[202]*(1)+in_buf[203]*(7)+in_buf[204]*(24)+in_buf[205]*(19)+in_buf[206]*(1)+in_buf[207]*(-15)+in_buf[208]*(-25)+in_buf[209]*(-14)+in_buf[210]*(9)+in_buf[211]*(12)+in_buf[212]*(4)+in_buf[213]*(9)+in_buf[214]*(12)+in_buf[215]*(10)+in_buf[216]*(14)+in_buf[217]*(21)+in_buf[218]*(18)+in_buf[219]*(-7)+in_buf[220]*(-9)+in_buf[221]*(5)+in_buf[222]*(25)+in_buf[223]*(8)+in_buf[224]*(-26)+in_buf[225]*(-18)+in_buf[226]*(17)+in_buf[227]*(7)+in_buf[228]*(-6)+in_buf[229]*(11)+in_buf[230]*(20)+in_buf[231]*(18)+in_buf[232]*(41)+in_buf[233]*(31)+in_buf[234]*(-4)+in_buf[235]*(-17)+in_buf[236]*(-22)+in_buf[237]*(-9)+in_buf[238]*(3)+in_buf[239]*(11)+in_buf[240]*(3)+in_buf[241]*(2)+in_buf[242]*(7)+in_buf[243]*(-4)+in_buf[244]*(3)+in_buf[245]*(10)+in_buf[246]*(-15)+in_buf[247]*(-22)+in_buf[248]*(15)+in_buf[249]*(30)+in_buf[250]*(28)+in_buf[251]*(-16)+in_buf[252]*(3)+in_buf[253]*(-9)+in_buf[254]*(-16)+in_buf[255]*(-5)+in_buf[256]*(6)+in_buf[257]*(5)+in_buf[258]*(16)+in_buf[259]*(22)+in_buf[260]*(33)+in_buf[261]*(23)+in_buf[262]*(-1)+in_buf[263]*(-6)+in_buf[264]*(-31)+in_buf[265]*(-31)+in_buf[266]*(-7)+in_buf[267]*(0)+in_buf[268]*(-1)+in_buf[269]*(-11)+in_buf[270]*(0)+in_buf[271]*(-3)+in_buf[272]*(10)+in_buf[273]*(7)+in_buf[274]*(-18)+in_buf[275]*(-12)+in_buf[276]*(10)+in_buf[277]*(20)+in_buf[278]*(15)+in_buf[279]*(-13)+in_buf[280]*(4)+in_buf[281]*(7)+in_buf[282]*(-30)+in_buf[283]*(-21)+in_buf[284]*(24)+in_buf[285]*(16)+in_buf[286]*(8)+in_buf[287]*(26)+in_buf[288]*(44)+in_buf[289]*(42)+in_buf[290]*(4)+in_buf[291]*(-16)+in_buf[292]*(-40)+in_buf[293]*(-47)+in_buf[294]*(-33)+in_buf[295]*(-7)+in_buf[296]*(-12)+in_buf[297]*(-16)+in_buf[298]*(-16)+in_buf[299]*(5)+in_buf[300]*(-15)+in_buf[301]*(-25)+in_buf[302]*(-21)+in_buf[303]*(-7)+in_buf[304]*(1)+in_buf[305]*(5)+in_buf[306]*(-24)+in_buf[307]*(-9)+in_buf[308]*(15)+in_buf[309]*(-9)+in_buf[310]*(-8)+in_buf[311]*(0)+in_buf[312]*(8)+in_buf[313]*(19)+in_buf[314]*(22)+in_buf[315]*(31)+in_buf[316]*(46)+in_buf[317]*(42)+in_buf[318]*(21)+in_buf[319]*(-3)+in_buf[320]*(-5)+in_buf[321]*(-23)+in_buf[322]*(-6)+in_buf[323]*(-1)+in_buf[324]*(-4)+in_buf[325]*(-27)+in_buf[326]*(-13)+in_buf[327]*(1)+in_buf[328]*(-15)+in_buf[329]*(-8)+in_buf[330]*(-18)+in_buf[331]*(-18)+in_buf[332]*(1)+in_buf[333]*(-2)+in_buf[334]*(-30)+in_buf[335]*(-28)+in_buf[336]*(26)+in_buf[337]*(15)+in_buf[338]*(-1)+in_buf[339]*(24)+in_buf[340]*(8)+in_buf[341]*(4)+in_buf[342]*(19)+in_buf[343]*(40)+in_buf[344]*(39)+in_buf[345]*(32)+in_buf[346]*(16)+in_buf[347]*(0)+in_buf[348]*(-18)+in_buf[349]*(-22)+in_buf[350]*(-12)+in_buf[351]*(5)+in_buf[352]*(0)+in_buf[353]*(-7)+in_buf[354]*(-6)+in_buf[355]*(-3)+in_buf[356]*(-8)+in_buf[357]*(3)+in_buf[358]*(-9)+in_buf[359]*(-16)+in_buf[360]*(13)+in_buf[361]*(-23)+in_buf[362]*(-37)+in_buf[363]*(-38)+in_buf[364]*(12)+in_buf[365]*(13)+in_buf[366]*(2)+in_buf[367]*(3)+in_buf[368]*(-9)+in_buf[369]*(11)+in_buf[370]*(13)+in_buf[371]*(35)+in_buf[372]*(36)+in_buf[373]*(23)+in_buf[374]*(13)+in_buf[375]*(-5)+in_buf[376]*(-20)+in_buf[377]*(-17)+in_buf[378]*(-1)+in_buf[379]*(8)+in_buf[380]*(-2)+in_buf[381]*(2)+in_buf[382]*(-1)+in_buf[383]*(0)+in_buf[384]*(0)+in_buf[385]*(1)+in_buf[386]*(9)+in_buf[387]*(3)+in_buf[388]*(-5)+in_buf[389]*(-35)+in_buf[390]*(-35)+in_buf[391]*(-16)+in_buf[392]*(13)+in_buf[393]*(10)+in_buf[394]*(17)+in_buf[395]*(-4)+in_buf[396]*(-2)+in_buf[397]*(23)+in_buf[398]*(20)+in_buf[399]*(24)+in_buf[400]*(28)+in_buf[401]*(23)+in_buf[402]*(7)+in_buf[403]*(-2)+in_buf[404]*(-21)+in_buf[405]*(-21)+in_buf[406]*(3)+in_buf[407]*(0)+in_buf[408]*(-4)+in_buf[409]*(2)+in_buf[410]*(-7)+in_buf[411]*(-5)+in_buf[412]*(-9)+in_buf[413]*(0)+in_buf[414]*(8)+in_buf[415]*(-7)+in_buf[416]*(-19)+in_buf[417]*(-28)+in_buf[418]*(-17)+in_buf[419]*(-11)+in_buf[420]*(10)+in_buf[421]*(2)+in_buf[422]*(26)+in_buf[423]*(25)+in_buf[424]*(2)+in_buf[425]*(5)+in_buf[426]*(21)+in_buf[427]*(26)+in_buf[428]*(28)+in_buf[429]*(14)+in_buf[430]*(6)+in_buf[431]*(-4)+in_buf[432]*(-8)+in_buf[433]*(-4)+in_buf[434]*(6)+in_buf[435]*(-3)+in_buf[436]*(3)+in_buf[437]*(-2)+in_buf[438]*(-13)+in_buf[439]*(-4)+in_buf[440]*(-8)+in_buf[441]*(-8)+in_buf[442]*(10)+in_buf[443]*(9)+in_buf[444]*(-41)+in_buf[445]*(0)+in_buf[446]*(3)+in_buf[447]*(-15)+in_buf[448]*(4)+in_buf[449]*(-2)+in_buf[450]*(7)+in_buf[451]*(27)+in_buf[452]*(1)+in_buf[453]*(10)+in_buf[454]*(22)+in_buf[455]*(7)+in_buf[456]*(15)+in_buf[457]*(2)+in_buf[458]*(-18)+in_buf[459]*(-26)+in_buf[460]*(-29)+in_buf[461]*(-10)+in_buf[462]*(8)+in_buf[463]*(14)+in_buf[464]*(27)+in_buf[465]*(-1)+in_buf[466]*(-12)+in_buf[467]*(5)+in_buf[468]*(9)+in_buf[469]*(2)+in_buf[470]*(7)+in_buf[471]*(2)+in_buf[472]*(-13)+in_buf[473]*(28)+in_buf[474]*(-30)+in_buf[475]*(-17)+in_buf[476]*(-2)+in_buf[477]*(-2)+in_buf[478]*(18)+in_buf[479]*(10)+in_buf[480]*(0)+in_buf[481]*(2)+in_buf[482]*(8)+in_buf[483]*(-14)+in_buf[484]*(3)+in_buf[485]*(-17)+in_buf[486]*(-13)+in_buf[487]*(-25)+in_buf[488]*(-20)+in_buf[489]*(10)+in_buf[490]*(29)+in_buf[491]*(29)+in_buf[492]*(26)+in_buf[493]*(8)+in_buf[494]*(3)+in_buf[495]*(7)+in_buf[496]*(21)+in_buf[497]*(-8)+in_buf[498]*(4)+in_buf[499]*(3)+in_buf[500]*(18)+in_buf[501]*(16)+in_buf[502]*(-14)+in_buf[503]*(-11)+in_buf[504]*(-31)+in_buf[505]*(-4)+in_buf[506]*(14)+in_buf[507]*(11)+in_buf[508]*(-1)+in_buf[509]*(1)+in_buf[510]*(5)+in_buf[511]*(-13)+in_buf[512]*(1)+in_buf[513]*(-6)+in_buf[514]*(-16)+in_buf[515]*(-24)+in_buf[516]*(-2)+in_buf[517]*(30)+in_buf[518]*(49)+in_buf[519]*(20)+in_buf[520]*(10)+in_buf[521]*(9)+in_buf[522]*(8)+in_buf[523]*(-5)+in_buf[524]*(4)+in_buf[525]*(-16)+in_buf[526]*(-11)+in_buf[527]*(-5)+in_buf[528]*(29)+in_buf[529]*(-4)+in_buf[530]*(-19)+in_buf[531]*(-3)+in_buf[532]*(0)+in_buf[533]*(-36)+in_buf[534]*(-24)+in_buf[535]*(-7)+in_buf[536]*(-29)+in_buf[537]*(-20)+in_buf[538]*(-4)+in_buf[539]*(-14)+in_buf[540]*(0)+in_buf[541]*(-3)+in_buf[542]*(-17)+in_buf[543]*(-7)+in_buf[544]*(7)+in_buf[545]*(26)+in_buf[546]*(40)+in_buf[547]*(20)+in_buf[548]*(4)+in_buf[549]*(1)+in_buf[550]*(11)+in_buf[551]*(-3)+in_buf[552]*(-3)+in_buf[553]*(-11)+in_buf[554]*(-10)+in_buf[555]*(8)+in_buf[556]*(36)+in_buf[557]*(2)+in_buf[558]*(-21)+in_buf[559]*(-5)+in_buf[560]*(1)+in_buf[561]*(0)+in_buf[562]*(1)+in_buf[563]*(-18)+in_buf[564]*(-44)+in_buf[565]*(-30)+in_buf[566]*(-8)+in_buf[567]*(-13)+in_buf[568]*(-10)+in_buf[569]*(-16)+in_buf[570]*(-8)+in_buf[571]*(1)+in_buf[572]*(35)+in_buf[573]*(15)+in_buf[574]*(19)+in_buf[575]*(20)+in_buf[576]*(6)+in_buf[577]*(11)+in_buf[578]*(24)+in_buf[579]*(-1)+in_buf[580]*(-14)+in_buf[581]*(-10)+in_buf[582]*(-9)+in_buf[583]*(-4)+in_buf[584]*(30)+in_buf[585]*(8)+in_buf[586]*(-15)+in_buf[587]*(4)+in_buf[588]*(-13)+in_buf[589]*(-5)+in_buf[590]*(-2)+in_buf[591]*(-4)+in_buf[592]*(-21)+in_buf[593]*(-19)+in_buf[594]*(-17)+in_buf[595]*(-4)+in_buf[596]*(7)+in_buf[597]*(0)+in_buf[598]*(-2)+in_buf[599]*(-2)+in_buf[600]*(16)+in_buf[601]*(17)+in_buf[602]*(20)+in_buf[603]*(20)+in_buf[604]*(9)+in_buf[605]*(32)+in_buf[606]*(9)+in_buf[607]*(-4)+in_buf[608]*(0)+in_buf[609]*(-3)+in_buf[610]*(-2)+in_buf[611]*(9)+in_buf[612]*(3)+in_buf[613]*(-2)+in_buf[614]*(-30)+in_buf[615]*(-3)+in_buf[616]*(-11)+in_buf[617]*(-13)+in_buf[618]*(-12)+in_buf[619]*(-20)+in_buf[620]*(4)+in_buf[621]*(-18)+in_buf[622]*(-26)+in_buf[623]*(-15)+in_buf[624]*(-13)+in_buf[625]*(-7)+in_buf[626]*(-1)+in_buf[627]*(-2)+in_buf[628]*(-7)+in_buf[629]*(0)+in_buf[630]*(13)+in_buf[631]*(17)+in_buf[632]*(8)+in_buf[633]*(12)+in_buf[634]*(4)+in_buf[635]*(10)+in_buf[636]*(-6)+in_buf[637]*(4)+in_buf[638]*(-3)+in_buf[639]*(20)+in_buf[640]*(17)+in_buf[641]*(0)+in_buf[642]*(10)+in_buf[643]*(-1)+in_buf[644]*(-3)+in_buf[645]*(3)+in_buf[646]*(0)+in_buf[647]*(-18)+in_buf[648]*(-20)+in_buf[649]*(-29)+in_buf[650]*(-38)+in_buf[651]*(-28)+in_buf[652]*(-14)+in_buf[653]*(-1)+in_buf[654]*(-4)+in_buf[655]*(-26)+in_buf[656]*(-7)+in_buf[657]*(-6)+in_buf[658]*(7)+in_buf[659]*(7)+in_buf[660]*(8)+in_buf[661]*(4)+in_buf[662]*(7)+in_buf[663]*(20)+in_buf[664]*(12)+in_buf[665]*(23)+in_buf[666]*(8)+in_buf[667]*(13)+in_buf[668]*(-12)+in_buf[669]*(-1)+in_buf[670]*(15)+in_buf[671]*(-3)+in_buf[672]*(4)+in_buf[673]*(-2)+in_buf[674]*(14)+in_buf[675]*(-13)+in_buf[676]*(-4)+in_buf[677]*(-19)+in_buf[678]*(-47)+in_buf[679]*(-33)+in_buf[680]*(-39)+in_buf[681]*(-5)+in_buf[682]*(-12)+in_buf[683]*(-13)+in_buf[684]*(-5)+in_buf[685]*(-13)+in_buf[686]*(-6)+in_buf[687]*(1)+in_buf[688]*(0)+in_buf[689]*(-15)+in_buf[690]*(11)+in_buf[691]*(35)+in_buf[692]*(22)+in_buf[693]*(18)+in_buf[694]*(27)+in_buf[695]*(6)+in_buf[696]*(-8)+in_buf[697]*(-3)+in_buf[698]*(-8)+in_buf[699]*(1)+in_buf[700]*(1)+in_buf[701]*(0)+in_buf[702]*(19)+in_buf[703]*(8)+in_buf[704]*(6)+in_buf[705]*(-23)+in_buf[706]*(-7)+in_buf[707]*(-20)+in_buf[708]*(-14)+in_buf[709]*(-11)+in_buf[710]*(-5)+in_buf[711]*(-8)+in_buf[712]*(-20)+in_buf[713]*(-5)+in_buf[714]*(11)+in_buf[715]*(18)+in_buf[716]*(0)+in_buf[717]*(20)+in_buf[718]*(35)+in_buf[719]*(8)+in_buf[720]*(18)+in_buf[721]*(51)+in_buf[722]*(45)+in_buf[723]*(11)+in_buf[724]*(-35)+in_buf[725]*(2)+in_buf[726]*(-4)+in_buf[727]*(0)+in_buf[728]*(-2)+in_buf[729]*(4)+in_buf[730]*(0)+in_buf[731]*(0)+in_buf[732]*(-10)+in_buf[733]*(-33)+in_buf[734]*(-28)+in_buf[735]*(-28)+in_buf[736]*(2)+in_buf[737]*(5)+in_buf[738]*(-39)+in_buf[739]*(-22)+in_buf[740]*(-1)+in_buf[741]*(13)+in_buf[742]*(4)+in_buf[743]*(11)+in_buf[744]*(-17)+in_buf[745]*(-12)+in_buf[746]*(-3)+in_buf[747]*(-21)+in_buf[748]*(-11)+in_buf[749]*(20)+in_buf[750]*(-4)+in_buf[751]*(11)+in_buf[752]*(-10)+in_buf[753]*(6)+in_buf[754]*(3)+in_buf[755]*(0)+in_buf[756]*(0)+in_buf[757]*(-1)+in_buf[758]*(0)+in_buf[759]*(4)+in_buf[760]*(14)+in_buf[761]*(18)+in_buf[762]*(7)+in_buf[763]*(-8)+in_buf[764]*(-13)+in_buf[765]*(13)+in_buf[766]*(-5)+in_buf[767]*(21)+in_buf[768]*(22)+in_buf[769]*(43)+in_buf[770]*(-16)+in_buf[771]*(-4)+in_buf[772]*(0)+in_buf[773]*(-9)+in_buf[774]*(-14)+in_buf[775]*(21)+in_buf[776]*(52)+in_buf[777]*(11)+in_buf[778]*(11)+in_buf[779]*(22)+in_buf[780]*(-2)+in_buf[781]*(4)+in_buf[782]*(0)+in_buf[783]*(3);
assign in_buf_weight042=in_buf[0]*(1)+in_buf[1]*(-3)+in_buf[2]*(1)+in_buf[3]*(4)+in_buf[4]*(2)+in_buf[5]*(-3)+in_buf[6]*(2)+in_buf[7]*(-2)+in_buf[8]*(-3)+in_buf[9]*(0)+in_buf[10]*(-2)+in_buf[11]*(0)+in_buf[12]*(1)+in_buf[13]*(-1)+in_buf[14]*(4)+in_buf[15]*(6)+in_buf[16]*(1)+in_buf[17]*(-3)+in_buf[18]*(2)+in_buf[19]*(1)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(-3)+in_buf[23]*(-3)+in_buf[24]*(1)+in_buf[25]*(-1)+in_buf[26]*(0)+in_buf[27]*(4)+in_buf[28]*(4)+in_buf[29]*(-3)+in_buf[30]*(4)+in_buf[31]*(-3)+in_buf[32]*(-3)+in_buf[33]*(3)+in_buf[34]*(2)+in_buf[35]*(0)+in_buf[36]*(0)+in_buf[37]*(-2)+in_buf[38]*(6)+in_buf[39]*(3)+in_buf[40]*(-6)+in_buf[41]*(-7)+in_buf[42]*(13)+in_buf[43]*(23)+in_buf[44]*(26)+in_buf[45]*(23)+in_buf[46]*(3)+in_buf[47]*(-5)+in_buf[48]*(-11)+in_buf[49]*(0)+in_buf[50]*(3)+in_buf[51]*(-1)+in_buf[52]*(3)+in_buf[53]*(4)+in_buf[54]*(0)+in_buf[55]*(5)+in_buf[56]*(4)+in_buf[57]*(0)+in_buf[58]*(-3)+in_buf[59]*(4)+in_buf[60]*(-2)+in_buf[61]*(1)+in_buf[62]*(1)+in_buf[63]*(-3)+in_buf[64]*(21)+in_buf[65]*(27)+in_buf[66]*(36)+in_buf[67]*(16)+in_buf[68]*(3)+in_buf[69]*(-11)+in_buf[70]*(-5)+in_buf[71]*(-20)+in_buf[72]*(-22)+in_buf[73]*(-3)+in_buf[74]*(-1)+in_buf[75]*(-38)+in_buf[76]*(-28)+in_buf[77]*(-30)+in_buf[78]*(-30)+in_buf[79]*(10)+in_buf[80]*(11)+in_buf[81]*(13)+in_buf[82]*(-1)+in_buf[83]*(1)+in_buf[84]*(0)+in_buf[85]*(-2)+in_buf[86]*(19)+in_buf[87]*(16)+in_buf[88]*(9)+in_buf[89]*(-6)+in_buf[90]*(6)+in_buf[91]*(25)+in_buf[92]*(40)+in_buf[93]*(57)+in_buf[94]*(40)+in_buf[95]*(27)+in_buf[96]*(32)+in_buf[97]*(-2)+in_buf[98]*(-29)+in_buf[99]*(-28)+in_buf[100]*(-13)+in_buf[101]*(-4)+in_buf[102]*(-11)+in_buf[103]*(-8)+in_buf[104]*(-11)+in_buf[105]*(-36)+in_buf[106]*(-21)+in_buf[107]*(2)+in_buf[108]*(38)+in_buf[109]*(35)+in_buf[110]*(20)+in_buf[111]*(4)+in_buf[112]*(0)+in_buf[113]*(-5)+in_buf[114]*(21)+in_buf[115]*(16)+in_buf[116]*(0)+in_buf[117]*(-7)+in_buf[118]*(19)+in_buf[119]*(9)+in_buf[120]*(3)+in_buf[121]*(9)+in_buf[122]*(-4)+in_buf[123]*(13)+in_buf[124]*(24)+in_buf[125]*(7)+in_buf[126]*(-5)+in_buf[127]*(-10)+in_buf[128]*(-23)+in_buf[129]*(-25)+in_buf[130]*(1)+in_buf[131]*(-9)+in_buf[132]*(0)+in_buf[133]*(-15)+in_buf[134]*(-13)+in_buf[135]*(5)+in_buf[136]*(-5)+in_buf[137]*(15)+in_buf[138]*(29)+in_buf[139]*(-14)+in_buf[140]*(-2)+in_buf[141]*(4)+in_buf[142]*(25)+in_buf[143]*(29)+in_buf[144]*(28)+in_buf[145]*(-7)+in_buf[146]*(-11)+in_buf[147]*(-15)+in_buf[148]*(2)+in_buf[149]*(0)+in_buf[150]*(4)+in_buf[151]*(7)+in_buf[152]*(0)+in_buf[153]*(15)+in_buf[154]*(7)+in_buf[155]*(-2)+in_buf[156]*(-1)+in_buf[157]*(-7)+in_buf[158]*(-10)+in_buf[159]*(-18)+in_buf[160]*(-5)+in_buf[161]*(-3)+in_buf[162]*(7)+in_buf[163]*(4)+in_buf[164]*(-3)+in_buf[165]*(31)+in_buf[166]*(-5)+in_buf[167]*(-18)+in_buf[168]*(3)+in_buf[169]*(10)+in_buf[170]*(0)+in_buf[171]*(31)+in_buf[172]*(17)+in_buf[173]*(-4)+in_buf[174]*(13)+in_buf[175]*(2)+in_buf[176]*(6)+in_buf[177]*(31)+in_buf[178]*(28)+in_buf[179]*(18)+in_buf[180]*(21)+in_buf[181]*(18)+in_buf[182]*(35)+in_buf[183]*(28)+in_buf[184]*(24)+in_buf[185]*(29)+in_buf[186]*(17)+in_buf[187]*(-7)+in_buf[188]*(3)+in_buf[189]*(10)+in_buf[190]*(-4)+in_buf[191]*(-5)+in_buf[192]*(18)+in_buf[193]*(28)+in_buf[194]*(-1)+in_buf[195]*(-16)+in_buf[196]*(1)+in_buf[197]*(6)+in_buf[198]*(25)+in_buf[199]*(56)+in_buf[200]*(19)+in_buf[201]*(-20)+in_buf[202]*(-1)+in_buf[203]*(0)+in_buf[204]*(21)+in_buf[205]*(10)+in_buf[206]*(24)+in_buf[207]*(18)+in_buf[208]*(30)+in_buf[209]*(32)+in_buf[210]*(53)+in_buf[211]*(40)+in_buf[212]*(42)+in_buf[213]*(30)+in_buf[214]*(30)+in_buf[215]*(7)+in_buf[216]*(15)+in_buf[217]*(14)+in_buf[218]*(6)+in_buf[219]*(-5)+in_buf[220]*(-8)+in_buf[221]*(12)+in_buf[222]*(15)+in_buf[223]*(-9)+in_buf[224]*(-16)+in_buf[225]*(8)+in_buf[226]*(8)+in_buf[227]*(2)+in_buf[228]*(2)+in_buf[229]*(-3)+in_buf[230]*(-12)+in_buf[231]*(1)+in_buf[232]*(21)+in_buf[233]*(10)+in_buf[234]*(20)+in_buf[235]*(17)+in_buf[236]*(28)+in_buf[237]*(34)+in_buf[238]*(57)+in_buf[239]*(49)+in_buf[240]*(33)+in_buf[241]*(26)+in_buf[242]*(25)+in_buf[243]*(5)+in_buf[244]*(3)+in_buf[245]*(-13)+in_buf[246]*(15)+in_buf[247]*(18)+in_buf[248]*(-2)+in_buf[249]*(28)+in_buf[250]*(37)+in_buf[251]*(25)+in_buf[252]*(12)+in_buf[253]*(10)+in_buf[254]*(10)+in_buf[255]*(10)+in_buf[256]*(10)+in_buf[257]*(0)+in_buf[258]*(6)+in_buf[259]*(7)+in_buf[260]*(11)+in_buf[261]*(4)+in_buf[262]*(14)+in_buf[263]*(6)+in_buf[264]*(24)+in_buf[265]*(34)+in_buf[266]*(35)+in_buf[267]*(28)+in_buf[268]*(12)+in_buf[269]*(8)+in_buf[270]*(0)+in_buf[271]*(0)+in_buf[272]*(-8)+in_buf[273]*(-23)+in_buf[274]*(0)+in_buf[275]*(20)+in_buf[276]*(20)+in_buf[277]*(52)+in_buf[278]*(58)+in_buf[279]*(27)+in_buf[280]*(16)+in_buf[281]*(10)+in_buf[282]*(21)+in_buf[283]*(13)+in_buf[284]*(-5)+in_buf[285]*(0)+in_buf[286]*(9)+in_buf[287]*(-3)+in_buf[288]*(14)+in_buf[289]*(0)+in_buf[290]*(-4)+in_buf[291]*(1)+in_buf[292]*(-7)+in_buf[293]*(0)+in_buf[294]*(-1)+in_buf[295]*(-12)+in_buf[296]*(0)+in_buf[297]*(-3)+in_buf[298]*(-3)+in_buf[299]*(-6)+in_buf[300]*(-4)+in_buf[301]*(-17)+in_buf[302]*(-24)+in_buf[303]*(-16)+in_buf[304]*(49)+in_buf[305]*(38)+in_buf[306]*(58)+in_buf[307]*(25)+in_buf[308]*(11)+in_buf[309]*(15)+in_buf[310]*(20)+in_buf[311]*(-2)+in_buf[312]*(-5)+in_buf[313]*(2)+in_buf[314]*(6)+in_buf[315]*(-12)+in_buf[316]*(-6)+in_buf[317]*(-20)+in_buf[318]*(-16)+in_buf[319]*(-7)+in_buf[320]*(-42)+in_buf[321]*(-47)+in_buf[322]*(-33)+in_buf[323]*(-22)+in_buf[324]*(-8)+in_buf[325]*(1)+in_buf[326]*(13)+in_buf[327]*(0)+in_buf[328]*(-2)+in_buf[329]*(-30)+in_buf[330]*(-27)+in_buf[331]*(4)+in_buf[332]*(3)+in_buf[333]*(6)+in_buf[334]*(39)+in_buf[335]*(0)+in_buf[336]*(0)+in_buf[337]*(0)+in_buf[338]*(14)+in_buf[339]*(-11)+in_buf[340]*(-13)+in_buf[341]*(-17)+in_buf[342]*(-19)+in_buf[343]*(-18)+in_buf[344]*(-13)+in_buf[345]*(-19)+in_buf[346]*(-28)+in_buf[347]*(-28)+in_buf[348]*(-54)+in_buf[349]*(-67)+in_buf[350]*(-22)+in_buf[351]*(-6)+in_buf[352]*(2)+in_buf[353]*(0)+in_buf[354]*(8)+in_buf[355]*(1)+in_buf[356]*(-4)+in_buf[357]*(-25)+in_buf[358]*(-46)+in_buf[359]*(-30)+in_buf[360]*(-18)+in_buf[361]*(-2)+in_buf[362]*(4)+in_buf[363]*(1)+in_buf[364]*(-21)+in_buf[365]*(13)+in_buf[366]*(24)+in_buf[367]*(-36)+in_buf[368]*(-41)+in_buf[369]*(-41)+in_buf[370]*(-20)+in_buf[371]*(-26)+in_buf[372]*(-19)+in_buf[373]*(-23)+in_buf[374]*(-28)+in_buf[375]*(-20)+in_buf[376]*(-32)+in_buf[377]*(-5)+in_buf[378]*(2)+in_buf[379]*(1)+in_buf[380]*(-1)+in_buf[381]*(6)+in_buf[382]*(3)+in_buf[383]*(1)+in_buf[384]*(-16)+in_buf[385]*(-16)+in_buf[386]*(-41)+in_buf[387]*(-39)+in_buf[388]*(-20)+in_buf[389]*(-15)+in_buf[390]*(4)+in_buf[391]*(7)+in_buf[392]*(-4)+in_buf[393]*(13)+in_buf[394]*(25)+in_buf[395]*(-33)+in_buf[396]*(-37)+in_buf[397]*(-54)+in_buf[398]*(-7)+in_buf[399]*(-18)+in_buf[400]*(-17)+in_buf[401]*(-23)+in_buf[402]*(-12)+in_buf[403]*(-20)+in_buf[404]*(-23)+in_buf[405]*(-2)+in_buf[406]*(10)+in_buf[407]*(10)+in_buf[408]*(-4)+in_buf[409]*(0)+in_buf[410]*(10)+in_buf[411]*(3)+in_buf[412]*(-18)+in_buf[413]*(-24)+in_buf[414]*(-30)+in_buf[415]*(-22)+in_buf[416]*(-16)+in_buf[417]*(-33)+in_buf[418]*(28)+in_buf[419]*(11)+in_buf[420]*(-3)+in_buf[421]*(-7)+in_buf[422]*(15)+in_buf[423]*(-31)+in_buf[424]*(-20)+in_buf[425]*(-40)+in_buf[426]*(-10)+in_buf[427]*(-10)+in_buf[428]*(-9)+in_buf[429]*(-19)+in_buf[430]*(-9)+in_buf[431]*(-10)+in_buf[432]*(-9)+in_buf[433]*(2)+in_buf[434]*(0)+in_buf[435]*(5)+in_buf[436]*(0)+in_buf[437]*(-1)+in_buf[438]*(8)+in_buf[439]*(-9)+in_buf[440]*(-17)+in_buf[441]*(-35)+in_buf[442]*(-33)+in_buf[443]*(-13)+in_buf[444]*(-1)+in_buf[445]*(-22)+in_buf[446]*(-2)+in_buf[447]*(24)+in_buf[448]*(4)+in_buf[449]*(-10)+in_buf[450]*(8)+in_buf[451]*(-10)+in_buf[452]*(-27)+in_buf[453]*(-38)+in_buf[454]*(-5)+in_buf[455]*(-12)+in_buf[456]*(-3)+in_buf[457]*(-10)+in_buf[458]*(2)+in_buf[459]*(10)+in_buf[460]*(2)+in_buf[461]*(13)+in_buf[462]*(-9)+in_buf[463]*(-12)+in_buf[464]*(-4)+in_buf[465]*(-10)+in_buf[466]*(-10)+in_buf[467]*(-16)+in_buf[468]*(-21)+in_buf[469]*(-10)+in_buf[470]*(-19)+in_buf[471]*(-21)+in_buf[472]*(-1)+in_buf[473]*(11)+in_buf[474]*(9)+in_buf[475]*(17)+in_buf[476]*(4)+in_buf[477]*(-7)+in_buf[478]*(2)+in_buf[479]*(0)+in_buf[480]*(-16)+in_buf[481]*(-12)+in_buf[482]*(0)+in_buf[483]*(-13)+in_buf[484]*(0)+in_buf[485]*(0)+in_buf[486]*(-7)+in_buf[487]*(-5)+in_buf[488]*(-6)+in_buf[489]*(5)+in_buf[490]*(1)+in_buf[491]*(3)+in_buf[492]*(3)+in_buf[493]*(-1)+in_buf[494]*(-2)+in_buf[495]*(-18)+in_buf[496]*(-16)+in_buf[497]*(-31)+in_buf[498]*(-33)+in_buf[499]*(-43)+in_buf[500]*(7)+in_buf[501]*(69)+in_buf[502]*(28)+in_buf[503]*(19)+in_buf[504]*(33)+in_buf[505]*(-5)+in_buf[506]*(5)+in_buf[507]*(4)+in_buf[508]*(5)+in_buf[509]*(8)+in_buf[510]*(20)+in_buf[511]*(11)+in_buf[512]*(7)+in_buf[513]*(-2)+in_buf[514]*(-11)+in_buf[515]*(-15)+in_buf[516]*(-6)+in_buf[517]*(2)+in_buf[518]*(6)+in_buf[519]*(10)+in_buf[520]*(3)+in_buf[521]*(9)+in_buf[522]*(2)+in_buf[523]*(-17)+in_buf[524]*(-15)+in_buf[525]*(-35)+in_buf[526]*(-16)+in_buf[527]*(-5)+in_buf[528]*(20)+in_buf[529]*(57)+in_buf[530]*(46)+in_buf[531]*(26)+in_buf[532]*(-18)+in_buf[533]*(4)+in_buf[534]*(2)+in_buf[535]*(-2)+in_buf[536]*(-5)+in_buf[537]*(1)+in_buf[538]*(30)+in_buf[539]*(20)+in_buf[540]*(18)+in_buf[541]*(2)+in_buf[542]*(2)+in_buf[543]*(-3)+in_buf[544]*(16)+in_buf[545]*(18)+in_buf[546]*(11)+in_buf[547]*(11)+in_buf[548]*(9)+in_buf[549]*(2)+in_buf[550]*(-4)+in_buf[551]*(1)+in_buf[552]*(-1)+in_buf[553]*(-25)+in_buf[554]*(-17)+in_buf[555]*(3)+in_buf[556]*(20)+in_buf[557]*(56)+in_buf[558]*(32)+in_buf[559]*(23)+in_buf[560]*(0)+in_buf[561]*(0)+in_buf[562]*(15)+in_buf[563]*(15)+in_buf[564]*(-4)+in_buf[565]*(20)+in_buf[566]*(24)+in_buf[567]*(16)+in_buf[568]*(35)+in_buf[569]*(20)+in_buf[570]*(17)+in_buf[571]*(19)+in_buf[572]*(13)+in_buf[573]*(13)+in_buf[574]*(0)+in_buf[575]*(11)+in_buf[576]*(13)+in_buf[577]*(7)+in_buf[578]*(4)+in_buf[579]*(7)+in_buf[580]*(13)+in_buf[581]*(-4)+in_buf[582]*(-17)+in_buf[583]*(8)+in_buf[584]*(24)+in_buf[585]*(51)+in_buf[586]*(10)+in_buf[587]*(1)+in_buf[588]*(6)+in_buf[589]*(11)+in_buf[590]*(29)+in_buf[591]*(21)+in_buf[592]*(14)+in_buf[593]*(16)+in_buf[594]*(0)+in_buf[595]*(-6)+in_buf[596]*(0)+in_buf[597]*(25)+in_buf[598]*(30)+in_buf[599]*(13)+in_buf[600]*(12)+in_buf[601]*(4)+in_buf[602]*(10)+in_buf[603]*(9)+in_buf[604]*(5)+in_buf[605]*(-4)+in_buf[606]*(9)+in_buf[607]*(19)+in_buf[608]*(20)+in_buf[609]*(5)+in_buf[610]*(1)+in_buf[611]*(22)+in_buf[612]*(59)+in_buf[613]*(45)+in_buf[614]*(31)+in_buf[615]*(0)+in_buf[616]*(8)+in_buf[617]*(-1)+in_buf[618]*(22)+in_buf[619]*(-5)+in_buf[620]*(21)+in_buf[621]*(36)+in_buf[622]*(7)+in_buf[623]*(-1)+in_buf[624]*(3)+in_buf[625]*(8)+in_buf[626]*(8)+in_buf[627]*(4)+in_buf[628]*(2)+in_buf[629]*(-6)+in_buf[630]*(7)+in_buf[631]*(-7)+in_buf[632]*(-4)+in_buf[633]*(-10)+in_buf[634]*(-10)+in_buf[635]*(-5)+in_buf[636]*(13)+in_buf[637]*(-4)+in_buf[638]*(2)+in_buf[639]*(36)+in_buf[640]*(62)+in_buf[641]*(32)+in_buf[642]*(7)+in_buf[643]*(-4)+in_buf[644]*(-2)+in_buf[645]*(-1)+in_buf[646]*(9)+in_buf[647]*(-22)+in_buf[648]*(16)+in_buf[649]*(24)+in_buf[650]*(25)+in_buf[651]*(5)+in_buf[652]*(-8)+in_buf[653]*(0)+in_buf[654]*(-7)+in_buf[655]*(7)+in_buf[656]*(0)+in_buf[657]*(-8)+in_buf[658]*(-10)+in_buf[659]*(-6)+in_buf[660]*(-6)+in_buf[661]*(-17)+in_buf[662]*(-23)+in_buf[663]*(-6)+in_buf[664]*(6)+in_buf[665]*(4)+in_buf[666]*(46)+in_buf[667]*(64)+in_buf[668]*(68)+in_buf[669]*(32)+in_buf[670]*(6)+in_buf[671]*(4)+in_buf[672]*(-2)+in_buf[673]*(0)+in_buf[674]*(14)+in_buf[675]*(11)+in_buf[676]*(33)+in_buf[677]*(18)+in_buf[678]*(-1)+in_buf[679]*(-9)+in_buf[680]*(-13)+in_buf[681]*(-8)+in_buf[682]*(-11)+in_buf[683]*(-3)+in_buf[684]*(12)+in_buf[685]*(4)+in_buf[686]*(-7)+in_buf[687]*(6)+in_buf[688]*(-16)+in_buf[689]*(-15)+in_buf[690]*(-13)+in_buf[691]*(5)+in_buf[692]*(17)+in_buf[693]*(20)+in_buf[694]*(6)+in_buf[695]*(23)+in_buf[696]*(49)+in_buf[697]*(0)+in_buf[698]*(4)+in_buf[699]*(-3)+in_buf[700]*(3)+in_buf[701]*(4)+in_buf[702]*(-32)+in_buf[703]*(30)+in_buf[704]*(25)+in_buf[705]*(7)+in_buf[706]*(-4)+in_buf[707]*(-10)+in_buf[708]*(33)+in_buf[709]*(36)+in_buf[710]*(12)+in_buf[711]*(16)+in_buf[712]*(31)+in_buf[713]*(26)+in_buf[714]*(32)+in_buf[715]*(20)+in_buf[716]*(19)+in_buf[717]*(21)+in_buf[718]*(18)+in_buf[719]*(19)+in_buf[720]*(16)+in_buf[721]*(25)+in_buf[722]*(14)+in_buf[723]*(34)+in_buf[724]*(42)+in_buf[725]*(0)+in_buf[726]*(11)+in_buf[727]*(0)+in_buf[728]*(-1)+in_buf[729]*(-1)+in_buf[730]*(4)+in_buf[731]*(16)+in_buf[732]*(-9)+in_buf[733]*(-29)+in_buf[734]*(-18)+in_buf[735]*(19)+in_buf[736]*(16)+in_buf[737]*(50)+in_buf[738]*(39)+in_buf[739]*(38)+in_buf[740]*(33)+in_buf[741]*(46)+in_buf[742]*(24)+in_buf[743]*(6)+in_buf[744]*(6)+in_buf[745]*(27)+in_buf[746]*(49)+in_buf[747]*(45)+in_buf[748]*(33)+in_buf[749]*(20)+in_buf[750]*(-1)+in_buf[751]*(13)+in_buf[752]*(3)+in_buf[753]*(14)+in_buf[754]*(-2)+in_buf[755]*(4)+in_buf[756]*(2)+in_buf[757]*(0)+in_buf[758]*(-1)+in_buf[759]*(-1)+in_buf[760]*(25)+in_buf[761]*(9)+in_buf[762]*(10)+in_buf[763]*(9)+in_buf[764]*(14)+in_buf[765]*(14)+in_buf[766]*(33)+in_buf[767]*(41)+in_buf[768]*(24)+in_buf[769]*(20)+in_buf[770]*(42)+in_buf[771]*(33)+in_buf[772]*(31)+in_buf[773]*(5)+in_buf[774]*(-11)+in_buf[775]*(-15)+in_buf[776]*(-1)+in_buf[777]*(-12)+in_buf[778]*(-16)+in_buf[779]*(6)+in_buf[780]*(2)+in_buf[781]*(-1)+in_buf[782]*(3)+in_buf[783]*(0);
assign in_buf_weight043=in_buf[0]*(3)+in_buf[1]*(0)+in_buf[2]*(1)+in_buf[3]*(0)+in_buf[4]*(1)+in_buf[5]*(4)+in_buf[6]*(-1)+in_buf[7]*(0)+in_buf[8]*(-4)+in_buf[9]*(-2)+in_buf[10]*(3)+in_buf[11]*(2)+in_buf[12]*(0)+in_buf[13]*(2)+in_buf[14]*(8)+in_buf[15]*(7)+in_buf[16]*(1)+in_buf[17]*(4)+in_buf[18]*(2)+in_buf[19]*(-2)+in_buf[20]*(4)+in_buf[21]*(1)+in_buf[22]*(-2)+in_buf[23]*(-3)+in_buf[24]*(3)+in_buf[25]*(-2)+in_buf[26]*(-2)+in_buf[27]*(0)+in_buf[28]*(-1)+in_buf[29]*(1)+in_buf[30]*(1)+in_buf[31]*(2)+in_buf[32]*(-1)+in_buf[33]*(2)+in_buf[34]*(0)+in_buf[35]*(-2)+in_buf[36]*(-3)+in_buf[37]*(1)+in_buf[38]*(-3)+in_buf[39]*(-2)+in_buf[40]*(-1)+in_buf[41]*(-2)+in_buf[42]*(-14)+in_buf[43]*(31)+in_buf[44]*(47)+in_buf[45]*(41)+in_buf[46]*(1)+in_buf[47]*(4)+in_buf[48]*(9)+in_buf[49]*(3)+in_buf[50]*(0)+in_buf[51]*(1)+in_buf[52]*(2)+in_buf[53]*(2)+in_buf[54]*(-3)+in_buf[55]*(4)+in_buf[56]*(2)+in_buf[57]*(-3)+in_buf[58]*(8)+in_buf[59]*(10)+in_buf[60]*(7)+in_buf[61]*(14)+in_buf[62]*(10)+in_buf[63]*(7)+in_buf[64]*(6)+in_buf[65]*(3)+in_buf[66]*(-13)+in_buf[67]*(-8)+in_buf[68]*(2)+in_buf[69]*(-9)+in_buf[70]*(10)+in_buf[71]*(39)+in_buf[72]*(57)+in_buf[73]*(42)+in_buf[74]*(14)+in_buf[75]*(-22)+in_buf[76]*(0)+in_buf[77]*(8)+in_buf[78]*(2)+in_buf[79]*(-12)+in_buf[80]*(-5)+in_buf[81]*(-7)+in_buf[82]*(4)+in_buf[83]*(-1)+in_buf[84]*(2)+in_buf[85]*(2)+in_buf[86]*(-14)+in_buf[87]*(6)+in_buf[88]*(6)+in_buf[89]*(7)+in_buf[90]*(8)+in_buf[91]*(-1)+in_buf[92]*(-16)+in_buf[93]*(-23)+in_buf[94]*(-48)+in_buf[95]*(-71)+in_buf[96]*(-56)+in_buf[97]*(-19)+in_buf[98]*(-10)+in_buf[99]*(6)+in_buf[100]*(5)+in_buf[101]*(11)+in_buf[102]*(22)+in_buf[103]*(-14)+in_buf[104]*(-20)+in_buf[105]*(17)+in_buf[106]*(14)+in_buf[107]*(32)+in_buf[108]*(20)+in_buf[109]*(-18)+in_buf[110]*(-34)+in_buf[111]*(-1)+in_buf[112]*(3)+in_buf[113]*(-5)+in_buf[114]*(-20)+in_buf[115]*(-15)+in_buf[116]*(-11)+in_buf[117]*(-8)+in_buf[118]*(-16)+in_buf[119]*(-37)+in_buf[120]*(-51)+in_buf[121]*(-40)+in_buf[122]*(-38)+in_buf[123]*(-35)+in_buf[124]*(-8)+in_buf[125]*(-5)+in_buf[126]*(11)+in_buf[127]*(18)+in_buf[128]*(29)+in_buf[129]*(22)+in_buf[130]*(-2)+in_buf[131]*(-5)+in_buf[132]*(3)+in_buf[133]*(7)+in_buf[134]*(-9)+in_buf[135]*(6)+in_buf[136]*(29)+in_buf[137]*(13)+in_buf[138]*(36)+in_buf[139]*(12)+in_buf[140]*(-3)+in_buf[141]*(0)+in_buf[142]*(6)+in_buf[143]*(-7)+in_buf[144]*(-7)+in_buf[145]*(-17)+in_buf[146]*(-32)+in_buf[147]*(-38)+in_buf[148]*(-53)+in_buf[149]*(-24)+in_buf[150]*(-14)+in_buf[151]*(10)+in_buf[152]*(11)+in_buf[153]*(9)+in_buf[154]*(10)+in_buf[155]*(4)+in_buf[156]*(6)+in_buf[157]*(19)+in_buf[158]*(15)+in_buf[159]*(16)+in_buf[160]*(27)+in_buf[161]*(16)+in_buf[162]*(1)+in_buf[163]*(-22)+in_buf[164]*(-1)+in_buf[165]*(24)+in_buf[166]*(32)+in_buf[167]*(1)+in_buf[168]*(1)+in_buf[169]*(-20)+in_buf[170]*(-1)+in_buf[171]*(-12)+in_buf[172]*(-24)+in_buf[173]*(-37)+in_buf[174]*(-68)+in_buf[175]*(-46)+in_buf[176]*(-35)+in_buf[177]*(-25)+in_buf[178]*(-14)+in_buf[179]*(8)+in_buf[180]*(8)+in_buf[181]*(6)+in_buf[182]*(6)+in_buf[183]*(11)+in_buf[184]*(11)+in_buf[185]*(20)+in_buf[186]*(9)+in_buf[187]*(14)+in_buf[188]*(7)+in_buf[189]*(-5)+in_buf[190]*(2)+in_buf[191]*(-9)+in_buf[192]*(-6)+in_buf[193]*(39)+in_buf[194]*(13)+in_buf[195]*(-16)+in_buf[196]*(0)+in_buf[197]*(-32)+in_buf[198]*(7)+in_buf[199]*(-20)+in_buf[200]*(-10)+in_buf[201]*(-33)+in_buf[202]*(-48)+in_buf[203]*(-52)+in_buf[204]*(-19)+in_buf[205]*(-10)+in_buf[206]*(0)+in_buf[207]*(7)+in_buf[208]*(7)+in_buf[209]*(3)+in_buf[210]*(-2)+in_buf[211]*(23)+in_buf[212]*(10)+in_buf[213]*(4)+in_buf[214]*(12)+in_buf[215]*(11)+in_buf[216]*(-2)+in_buf[217]*(13)+in_buf[218]*(8)+in_buf[219]*(-3)+in_buf[220]*(8)+in_buf[221]*(41)+in_buf[222]*(-4)+in_buf[223]*(-24)+in_buf[224]*(13)+in_buf[225]*(-18)+in_buf[226]*(-4)+in_buf[227]*(-8)+in_buf[228]*(-14)+in_buf[229]*(-39)+in_buf[230]*(-15)+in_buf[231]*(-24)+in_buf[232]*(-6)+in_buf[233]*(-3)+in_buf[234]*(5)+in_buf[235]*(19)+in_buf[236]*(1)+in_buf[237]*(5)+in_buf[238]*(-6)+in_buf[239]*(1)+in_buf[240]*(2)+in_buf[241]*(-5)+in_buf[242]*(1)+in_buf[243]*(12)+in_buf[244]*(1)+in_buf[245]*(12)+in_buf[246]*(0)+in_buf[247]*(10)+in_buf[248]*(28)+in_buf[249]*(34)+in_buf[250]*(16)+in_buf[251]*(11)+in_buf[252]*(0)+in_buf[253]*(-24)+in_buf[254]*(-15)+in_buf[255]*(-17)+in_buf[256]*(-41)+in_buf[257]*(-54)+in_buf[258]*(-18)+in_buf[259]*(-17)+in_buf[260]*(-7)+in_buf[261]*(12)+in_buf[262]*(21)+in_buf[263]*(15)+in_buf[264]*(2)+in_buf[265]*(12)+in_buf[266]*(-8)+in_buf[267]*(-15)+in_buf[268]*(-15)+in_buf[269]*(-18)+in_buf[270]*(-24)+in_buf[271]*(-1)+in_buf[272]*(1)+in_buf[273]*(0)+in_buf[274]*(-3)+in_buf[275]*(7)+in_buf[276]*(30)+in_buf[277]*(31)+in_buf[278]*(5)+in_buf[279]*(-18)+in_buf[280]*(1)+in_buf[281]*(-14)+in_buf[282]*(-31)+in_buf[283]*(-49)+in_buf[284]*(-41)+in_buf[285]*(-48)+in_buf[286]*(-5)+in_buf[287]*(-2)+in_buf[288]*(5)+in_buf[289]*(13)+in_buf[290]*(13)+in_buf[291]*(12)+in_buf[292]*(17)+in_buf[293]*(-2)+in_buf[294]*(-7)+in_buf[295]*(-20)+in_buf[296]*(-25)+in_buf[297]*(-29)+in_buf[298]*(-15)+in_buf[299]*(-6)+in_buf[300]*(0)+in_buf[301]*(-4)+in_buf[302]*(0)+in_buf[303]*(34)+in_buf[304]*(16)+in_buf[305]*(-10)+in_buf[306]*(8)+in_buf[307]*(0)+in_buf[308]*(0)+in_buf[309]*(-20)+in_buf[310]*(-29)+in_buf[311]*(-62)+in_buf[312]*(-46)+in_buf[313]*(-11)+in_buf[314]*(16)+in_buf[315]*(15)+in_buf[316]*(10)+in_buf[317]*(4)+in_buf[318]*(2)+in_buf[319]*(4)+in_buf[320]*(10)+in_buf[321]*(11)+in_buf[322]*(5)+in_buf[323]*(-13)+in_buf[324]*(-10)+in_buf[325]*(-10)+in_buf[326]*(-3)+in_buf[327]*(4)+in_buf[328]*(2)+in_buf[329]*(4)+in_buf[330]*(-4)+in_buf[331]*(21)+in_buf[332]*(36)+in_buf[333]*(30)+in_buf[334]*(41)+in_buf[335]*(-30)+in_buf[336]*(-5)+in_buf[337]*(-6)+in_buf[338]*(-4)+in_buf[339]*(-46)+in_buf[340]*(-29)+in_buf[341]*(-4)+in_buf[342]*(13)+in_buf[343]*(7)+in_buf[344]*(0)+in_buf[345]*(12)+in_buf[346]*(-6)+in_buf[347]*(5)+in_buf[348]*(1)+in_buf[349]*(17)+in_buf[350]*(11)+in_buf[351]*(2)+in_buf[352]*(0)+in_buf[353]*(15)+in_buf[354]*(5)+in_buf[355]*(22)+in_buf[356]*(21)+in_buf[357]*(17)+in_buf[358]*(-5)+in_buf[359]*(11)+in_buf[360]*(14)+in_buf[361]*(-6)+in_buf[362]*(8)+in_buf[363]*(-34)+in_buf[364]*(19)+in_buf[365]*(-7)+in_buf[366]*(-36)+in_buf[367]*(-46)+in_buf[368]*(-36)+in_buf[369]*(-21)+in_buf[370]*(-5)+in_buf[371]*(-1)+in_buf[372]*(-4)+in_buf[373]*(8)+in_buf[374]*(-2)+in_buf[375]*(9)+in_buf[376]*(21)+in_buf[377]*(24)+in_buf[378]*(22)+in_buf[379]*(24)+in_buf[380]*(11)+in_buf[381]*(1)+in_buf[382]*(1)+in_buf[383]*(12)+in_buf[384]*(-1)+in_buf[385]*(-13)+in_buf[386]*(1)+in_buf[387]*(-10)+in_buf[388]*(-36)+in_buf[389]*(-1)+in_buf[390]*(26)+in_buf[391]*(16)+in_buf[392]*(9)+in_buf[393]*(-15)+in_buf[394]*(-26)+in_buf[395]*(-40)+in_buf[396]*(-29)+in_buf[397]*(-12)+in_buf[398]*(-1)+in_buf[399]*(-7)+in_buf[400]*(-8)+in_buf[401]*(-4)+in_buf[402]*(1)+in_buf[403]*(18)+in_buf[404]*(16)+in_buf[405]*(25)+in_buf[406]*(13)+in_buf[407]*(12)+in_buf[408]*(13)+in_buf[409]*(6)+in_buf[410]*(-5)+in_buf[411]*(-24)+in_buf[412]*(-29)+in_buf[413]*(-18)+in_buf[414]*(-31)+in_buf[415]*(-35)+in_buf[416]*(-26)+in_buf[417]*(24)+in_buf[418]*(45)+in_buf[419]*(13)+in_buf[420]*(2)+in_buf[421]*(-8)+in_buf[422]*(-32)+in_buf[423]*(-40)+in_buf[424]*(-20)+in_buf[425]*(2)+in_buf[426]*(3)+in_buf[427]*(-4)+in_buf[428]*(-4)+in_buf[429]*(0)+in_buf[430]*(11)+in_buf[431]*(19)+in_buf[432]*(12)+in_buf[433]*(17)+in_buf[434]*(12)+in_buf[435]*(3)+in_buf[436]*(9)+in_buf[437]*(0)+in_buf[438]*(-8)+in_buf[439]*(-21)+in_buf[440]*(-36)+in_buf[441]*(-37)+in_buf[442]*(-25)+in_buf[443]*(-29)+in_buf[444]*(2)+in_buf[445]*(35)+in_buf[446]*(7)+in_buf[447]*(19)+in_buf[448]*(-6)+in_buf[449]*(-11)+in_buf[450]*(-39)+in_buf[451]*(-33)+in_buf[452]*(-33)+in_buf[453]*(-19)+in_buf[454]*(-2)+in_buf[455]*(-7)+in_buf[456]*(11)+in_buf[457]*(2)+in_buf[458]*(21)+in_buf[459]*(22)+in_buf[460]*(19)+in_buf[461]*(10)+in_buf[462]*(8)+in_buf[463]*(2)+in_buf[464]*(13)+in_buf[465]*(2)+in_buf[466]*(-10)+in_buf[467]*(-34)+in_buf[468]*(-39)+in_buf[469]*(-25)+in_buf[470]*(-5)+in_buf[471]*(-4)+in_buf[472]*(-2)+in_buf[473]*(62)+in_buf[474]*(41)+in_buf[475]*(11)+in_buf[476]*(-2)+in_buf[477]*(-9)+in_buf[478]*(-40)+in_buf[479]*(-22)+in_buf[480]*(-7)+in_buf[481]*(-6)+in_buf[482]*(-3)+in_buf[483]*(-3)+in_buf[484]*(10)+in_buf[485]*(19)+in_buf[486]*(18)+in_buf[487]*(16)+in_buf[488]*(14)+in_buf[489]*(-1)+in_buf[490]*(-2)+in_buf[491]*(3)+in_buf[492]*(7)+in_buf[493]*(4)+in_buf[494]*(-17)+in_buf[495]*(-34)+in_buf[496]*(-21)+in_buf[497]*(-24)+in_buf[498]*(-5)+in_buf[499]*(0)+in_buf[500]*(19)+in_buf[501]*(-3)+in_buf[502]*(17)+in_buf[503]*(27)+in_buf[504]*(22)+in_buf[505]*(-7)+in_buf[506]*(-43)+in_buf[507]*(-19)+in_buf[508]*(11)+in_buf[509]*(15)+in_buf[510]*(16)+in_buf[511]*(11)+in_buf[512]*(13)+in_buf[513]*(16)+in_buf[514]*(16)+in_buf[515]*(-3)+in_buf[516]*(-2)+in_buf[517]*(-11)+in_buf[518]*(-9)+in_buf[519]*(-2)+in_buf[520]*(-8)+in_buf[521]*(-2)+in_buf[522]*(-25)+in_buf[523]*(-20)+in_buf[524]*(-13)+in_buf[525]*(-29)+in_buf[526]*(-3)+in_buf[527]*(7)+in_buf[528]*(22)+in_buf[529]*(-12)+in_buf[530]*(-15)+in_buf[531]*(4)+in_buf[532]*(-5)+in_buf[533]*(-31)+in_buf[534]*(-13)+in_buf[535]*(-25)+in_buf[536]*(0)+in_buf[537]*(10)+in_buf[538]*(0)+in_buf[539]*(-1)+in_buf[540]*(13)+in_buf[541]*(2)+in_buf[542]*(0)+in_buf[543]*(-19)+in_buf[544]*(-25)+in_buf[545]*(-22)+in_buf[546]*(-24)+in_buf[547]*(3)+in_buf[548]*(4)+in_buf[549]*(2)+in_buf[550]*(7)+in_buf[551]*(0)+in_buf[552]*(-3)+in_buf[553]*(-15)+in_buf[554]*(14)+in_buf[555]*(32)+in_buf[556]*(23)+in_buf[557]*(-9)+in_buf[558]*(23)+in_buf[559]*(0)+in_buf[560]*(3)+in_buf[561]*(19)+in_buf[562]*(12)+in_buf[563]*(-9)+in_buf[564]*(0)+in_buf[565]*(12)+in_buf[566]*(5)+in_buf[567]*(7)+in_buf[568]*(14)+in_buf[569]*(0)+in_buf[570]*(0)+in_buf[571]*(-12)+in_buf[572]*(-24)+in_buf[573]*(-20)+in_buf[574]*(-25)+in_buf[575]*(0)+in_buf[576]*(-3)+in_buf[577]*(3)+in_buf[578]*(-1)+in_buf[579]*(-1)+in_buf[580]*(3)+in_buf[581]*(4)+in_buf[582]*(21)+in_buf[583]*(23)+in_buf[584]*(17)+in_buf[585]*(29)+in_buf[586]*(9)+in_buf[587]*(7)+in_buf[588]*(-26)+in_buf[589]*(-3)+in_buf[590]*(-17)+in_buf[591]*(-4)+in_buf[592]*(15)+in_buf[593]*(12)+in_buf[594]*(23)+in_buf[595]*(20)+in_buf[596]*(0)+in_buf[597]*(4)+in_buf[598]*(-7)+in_buf[599]*(-9)+in_buf[600]*(-16)+in_buf[601]*(-7)+in_buf[602]*(-14)+in_buf[603]*(-5)+in_buf[604]*(-7)+in_buf[605]*(18)+in_buf[606]*(-7)+in_buf[607]*(-1)+in_buf[608]*(-8)+in_buf[609]*(-13)+in_buf[610]*(13)+in_buf[611]*(11)+in_buf[612]*(-6)+in_buf[613]*(16)+in_buf[614]*(30)+in_buf[615]*(-5)+in_buf[616]*(-23)+in_buf[617]*(-12)+in_buf[618]*(-17)+in_buf[619]*(14)+in_buf[620]*(21)+in_buf[621]*(-2)+in_buf[622]*(18)+in_buf[623]*(18)+in_buf[624]*(1)+in_buf[625]*(5)+in_buf[626]*(0)+in_buf[627]*(13)+in_buf[628]*(11)+in_buf[629]*(19)+in_buf[630]*(6)+in_buf[631]*(0)+in_buf[632]*(9)+in_buf[633]*(2)+in_buf[634]*(-8)+in_buf[635]*(-15)+in_buf[636]*(-19)+in_buf[637]*(-24)+in_buf[638]*(-17)+in_buf[639]*(10)+in_buf[640]*(10)+in_buf[641]*(20)+in_buf[642]*(-1)+in_buf[643]*(-3)+in_buf[644]*(0)+in_buf[645]*(-3)+in_buf[646]*(-22)+in_buf[647]*(35)+in_buf[648]*(13)+in_buf[649]*(-5)+in_buf[650]*(-8)+in_buf[651]*(-13)+in_buf[652]*(7)+in_buf[653]*(-2)+in_buf[654]*(-3)+in_buf[655]*(2)+in_buf[656]*(15)+in_buf[657]*(19)+in_buf[658]*(10)+in_buf[659]*(21)+in_buf[660]*(17)+in_buf[661]*(3)+in_buf[662]*(0)+in_buf[663]*(-15)+in_buf[664]*(-21)+in_buf[665]*(-25)+in_buf[666]*(2)+in_buf[667]*(35)+in_buf[668]*(15)+in_buf[669]*(17)+in_buf[670]*(-14)+in_buf[671]*(3)+in_buf[672]*(3)+in_buf[673]*(-1)+in_buf[674]*(-1)+in_buf[675]*(-10)+in_buf[676]*(-19)+in_buf[677]*(-11)+in_buf[678]*(-9)+in_buf[679]*(-10)+in_buf[680]*(-8)+in_buf[681]*(-5)+in_buf[682]*(6)+in_buf[683]*(5)+in_buf[684]*(21)+in_buf[685]*(12)+in_buf[686]*(0)+in_buf[687]*(24)+in_buf[688]*(24)+in_buf[689]*(2)+in_buf[690]*(11)+in_buf[691]*(9)+in_buf[692]*(12)+in_buf[693]*(-12)+in_buf[694]*(-7)+in_buf[695]*(0)+in_buf[696]*(18)+in_buf[697]*(-4)+in_buf[698]*(-12)+in_buf[699]*(4)+in_buf[700]*(3)+in_buf[701]*(0)+in_buf[702]*(26)+in_buf[703]*(-11)+in_buf[704]*(-43)+in_buf[705]*(-27)+in_buf[706]*(-7)+in_buf[707]*(0)+in_buf[708]*(-8)+in_buf[709]*(1)+in_buf[710]*(10)+in_buf[711]*(-4)+in_buf[712]*(-5)+in_buf[713]*(6)+in_buf[714]*(14)+in_buf[715]*(21)+in_buf[716]*(36)+in_buf[717]*(54)+in_buf[718]*(40)+in_buf[719]*(54)+in_buf[720]*(41)+in_buf[721]*(23)+in_buf[722]*(-6)+in_buf[723]*(-23)+in_buf[724]*(-5)+in_buf[725]*(9)+in_buf[726]*(-10)+in_buf[727]*(2)+in_buf[728]*(1)+in_buf[729]*(-2)+in_buf[730]*(4)+in_buf[731]*(18)+in_buf[732]*(24)+in_buf[733]*(24)+in_buf[734]*(3)+in_buf[735]*(14)+in_buf[736]*(23)+in_buf[737]*(12)+in_buf[738]*(16)+in_buf[739]*(21)+in_buf[740]*(18)+in_buf[741]*(0)+in_buf[742]*(33)+in_buf[743]*(15)+in_buf[744]*(23)+in_buf[745]*(46)+in_buf[746]*(41)+in_buf[747]*(9)+in_buf[748]*(35)+in_buf[749]*(9)+in_buf[750]*(0)+in_buf[751]*(14)+in_buf[752]*(19)+in_buf[753]*(-4)+in_buf[754]*(3)+in_buf[755]*(-2)+in_buf[756]*(1)+in_buf[757]*(-1)+in_buf[758]*(4)+in_buf[759]*(-3)+in_buf[760]*(-19)+in_buf[761]*(-19)+in_buf[762]*(6)+in_buf[763]*(16)+in_buf[764]*(6)+in_buf[765]*(-6)+in_buf[766]*(-7)+in_buf[767]*(16)+in_buf[768]*(11)+in_buf[769]*(-2)+in_buf[770]*(29)+in_buf[771]*(21)+in_buf[772]*(4)+in_buf[773]*(19)+in_buf[774]*(39)+in_buf[775]*(25)+in_buf[776]*(7)+in_buf[777]*(-12)+in_buf[778]*(-15)+in_buf[779]*(-3)+in_buf[780]*(4)+in_buf[781]*(4)+in_buf[782]*(-3)+in_buf[783]*(4);
assign in_buf_weight044=in_buf[0]*(3)+in_buf[1]*(-1)+in_buf[2]*(4)+in_buf[3]*(0)+in_buf[4]*(4)+in_buf[5]*(3)+in_buf[6]*(1)+in_buf[7]*(-2)+in_buf[8]*(-2)+in_buf[9]*(1)+in_buf[10]*(3)+in_buf[11]*(0)+in_buf[12]*(7)+in_buf[13]*(3)+in_buf[14]*(-5)+in_buf[15]*(-1)+in_buf[16]*(-1)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(0)+in_buf[22]*(-1)+in_buf[23]*(-2)+in_buf[24]*(5)+in_buf[25]*(2)+in_buf[26]*(1)+in_buf[27]*(1)+in_buf[28]*(0)+in_buf[29]*(0)+in_buf[30]*(-1)+in_buf[31]*(1)+in_buf[32]*(8)+in_buf[33]*(2)+in_buf[34]*(4)+in_buf[35]*(8)+in_buf[36]*(10)+in_buf[37]*(3)+in_buf[38]*(6)+in_buf[39]*(1)+in_buf[40]*(10)+in_buf[41]*(13)+in_buf[42]*(27)+in_buf[43]*(12)+in_buf[44]*(3)+in_buf[45]*(9)+in_buf[46]*(37)+in_buf[47]*(19)+in_buf[48]*(18)+in_buf[49]*(8)+in_buf[50]*(10)+in_buf[51]*(7)+in_buf[52]*(0)+in_buf[53]*(0)+in_buf[54]*(-2)+in_buf[55]*(-3)+in_buf[56]*(-2)+in_buf[57]*(1)+in_buf[58]*(14)+in_buf[59]*(5)+in_buf[60]*(12)+in_buf[61]*(17)+in_buf[62]*(11)+in_buf[63]*(15)+in_buf[64]*(18)+in_buf[65]*(44)+in_buf[66]*(35)+in_buf[67]*(33)+in_buf[68]*(53)+in_buf[69]*(60)+in_buf[70]*(69)+in_buf[71]*(75)+in_buf[72]*(58)+in_buf[73]*(13)+in_buf[74]*(-12)+in_buf[75]*(4)+in_buf[76]*(-6)+in_buf[77]*(2)+in_buf[78]*(9)+in_buf[79]*(5)+in_buf[80]*(7)+in_buf[81]*(-1)+in_buf[82]*(0)+in_buf[83]*(-1)+in_buf[84]*(0)+in_buf[85]*(1)+in_buf[86]*(19)+in_buf[87]*(11)+in_buf[88]*(2)+in_buf[89]*(1)+in_buf[90]*(-12)+in_buf[91]*(-23)+in_buf[92]*(-27)+in_buf[93]*(5)+in_buf[94]*(5)+in_buf[95]*(1)+in_buf[96]*(-8)+in_buf[97]*(-12)+in_buf[98]*(-15)+in_buf[99]*(-9)+in_buf[100]*(13)+in_buf[101]*(8)+in_buf[102]*(1)+in_buf[103]*(45)+in_buf[104]*(18)+in_buf[105]*(5)+in_buf[106]*(29)+in_buf[107]*(33)+in_buf[108]*(5)+in_buf[109]*(-28)+in_buf[110]*(-9)+in_buf[111]*(-3)+in_buf[112]*(0)+in_buf[113]*(1)+in_buf[114]*(12)+in_buf[115]*(-33)+in_buf[116]*(-28)+in_buf[117]*(-32)+in_buf[118]*(-31)+in_buf[119]*(-25)+in_buf[120]*(-3)+in_buf[121]*(3)+in_buf[122]*(0)+in_buf[123]*(-13)+in_buf[124]*(0)+in_buf[125]*(1)+in_buf[126]*(1)+in_buf[127]*(0)+in_buf[128]*(5)+in_buf[129]*(16)+in_buf[130]*(0)+in_buf[131]*(16)+in_buf[132]*(12)+in_buf[133]*(6)+in_buf[134]*(13)+in_buf[135]*(-6)+in_buf[136]*(-30)+in_buf[137]*(-56)+in_buf[138]*(-19)+in_buf[139]*(2)+in_buf[140]*(-3)+in_buf[141]*(0)+in_buf[142]*(26)+in_buf[143]*(-11)+in_buf[144]*(-23)+in_buf[145]*(-30)+in_buf[146]*(-23)+in_buf[147]*(1)+in_buf[148]*(16)+in_buf[149]*(-2)+in_buf[150]*(-16)+in_buf[151]*(-5)+in_buf[152]*(16)+in_buf[153]*(8)+in_buf[154]*(0)+in_buf[155]*(11)+in_buf[156]*(2)+in_buf[157]*(5)+in_buf[158]*(1)+in_buf[159]*(-4)+in_buf[160]*(-13)+in_buf[161]*(11)+in_buf[162]*(9)+in_buf[163]*(6)+in_buf[164]*(8)+in_buf[165]*(-8)+in_buf[166]*(-1)+in_buf[167]*(6)+in_buf[168]*(1)+in_buf[169]*(0)+in_buf[170]*(-1)+in_buf[171]*(-8)+in_buf[172]*(-23)+in_buf[173]*(-34)+in_buf[174]*(-16)+in_buf[175]*(7)+in_buf[176]*(-22)+in_buf[177]*(-11)+in_buf[178]*(-19)+in_buf[179]*(-9)+in_buf[180]*(8)+in_buf[181]*(1)+in_buf[182]*(1)+in_buf[183]*(-4)+in_buf[184]*(-12)+in_buf[185]*(-13)+in_buf[186]*(-14)+in_buf[187]*(-11)+in_buf[188]*(-13)+in_buf[189]*(6)+in_buf[190]*(16)+in_buf[191]*(7)+in_buf[192]*(-12)+in_buf[193]*(-2)+in_buf[194]*(13)+in_buf[195]*(29)+in_buf[196]*(4)+in_buf[197]*(22)+in_buf[198]*(-9)+in_buf[199]*(-8)+in_buf[200]*(-13)+in_buf[201]*(2)+in_buf[202]*(-5)+in_buf[203]*(-18)+in_buf[204]*(-30)+in_buf[205]*(-14)+in_buf[206]*(-12)+in_buf[207]*(-6)+in_buf[208]*(-3)+in_buf[209]*(6)+in_buf[210]*(-1)+in_buf[211]*(-5)+in_buf[212]*(-6)+in_buf[213]*(-3)+in_buf[214]*(0)+in_buf[215]*(-2)+in_buf[216]*(-2)+in_buf[217]*(10)+in_buf[218]*(29)+in_buf[219]*(9)+in_buf[220]*(-15)+in_buf[221]*(-33)+in_buf[222]*(-4)+in_buf[223]*(20)+in_buf[224]*(1)+in_buf[225]*(20)+in_buf[226]*(-13)+in_buf[227]*(-7)+in_buf[228]*(-6)+in_buf[229]*(15)+in_buf[230]*(11)+in_buf[231]*(0)+in_buf[232]*(1)+in_buf[233]*(-1)+in_buf[234]*(-5)+in_buf[235]*(0)+in_buf[236]*(12)+in_buf[237]*(22)+in_buf[238]*(9)+in_buf[239]*(5)+in_buf[240]*(-17)+in_buf[241]*(0)+in_buf[242]*(-16)+in_buf[243]*(-3)+in_buf[244]*(-9)+in_buf[245]*(0)+in_buf[246]*(17)+in_buf[247]*(9)+in_buf[248]*(-34)+in_buf[249]*(-29)+in_buf[250]*(8)+in_buf[251]*(-24)+in_buf[252]*(4)+in_buf[253]*(14)+in_buf[254]*(-3)+in_buf[255]*(14)+in_buf[256]*(-12)+in_buf[257]*(-10)+in_buf[258]*(-2)+in_buf[259]*(-6)+in_buf[260]*(3)+in_buf[261]*(15)+in_buf[262]*(-1)+in_buf[263]*(0)+in_buf[264]*(6)+in_buf[265]*(1)+in_buf[266]*(4)+in_buf[267]*(9)+in_buf[268]*(-7)+in_buf[269]*(-11)+in_buf[270]*(-6)+in_buf[271]*(-15)+in_buf[272]*(-18)+in_buf[273]*(-3)+in_buf[274]*(1)+in_buf[275]*(1)+in_buf[276]*(-9)+in_buf[277]*(10)+in_buf[278]*(5)+in_buf[279]*(27)+in_buf[280]*(0)+in_buf[281]*(11)+in_buf[282]*(-11)+in_buf[283]*(-7)+in_buf[284]*(-28)+in_buf[285]*(-19)+in_buf[286]*(-9)+in_buf[287]*(-8)+in_buf[288]*(5)+in_buf[289]*(11)+in_buf[290]*(0)+in_buf[291]*(2)+in_buf[292]*(0)+in_buf[293]*(9)+in_buf[294]*(9)+in_buf[295]*(5)+in_buf[296]*(-5)+in_buf[297]*(-9)+in_buf[298]*(-6)+in_buf[299]*(-3)+in_buf[300]*(-17)+in_buf[301]*(-4)+in_buf[302]*(-20)+in_buf[303]*(-14)+in_buf[304]*(9)+in_buf[305]*(-4)+in_buf[306]*(-1)+in_buf[307]*(31)+in_buf[308]*(-1)+in_buf[309]*(6)+in_buf[310]*(1)+in_buf[311]*(-26)+in_buf[312]*(-13)+in_buf[313]*(-4)+in_buf[314]*(-2)+in_buf[315]*(1)+in_buf[316]*(15)+in_buf[317]*(23)+in_buf[318]*(-3)+in_buf[319]*(2)+in_buf[320]*(3)+in_buf[321]*(19)+in_buf[322]*(22)+in_buf[323]*(10)+in_buf[324]*(-7)+in_buf[325]*(-28)+in_buf[326]*(-25)+in_buf[327]*(-19)+in_buf[328]*(0)+in_buf[329]*(-4)+in_buf[330]*(-15)+in_buf[331]*(8)+in_buf[332]*(-5)+in_buf[333]*(-22)+in_buf[334]*(-34)+in_buf[335]*(34)+in_buf[336]*(1)+in_buf[337]*(1)+in_buf[338]*(11)+in_buf[339]*(-21)+in_buf[340]*(6)+in_buf[341]*(-17)+in_buf[342]*(-18)+in_buf[343]*(-16)+in_buf[344]*(16)+in_buf[345]*(15)+in_buf[346]*(-15)+in_buf[347]*(-1)+in_buf[348]*(11)+in_buf[349]*(4)+in_buf[350]*(18)+in_buf[351]*(18)+in_buf[352]*(3)+in_buf[353]*(-12)+in_buf[354]*(-15)+in_buf[355]*(-18)+in_buf[356]*(2)+in_buf[357]*(-8)+in_buf[358]*(12)+in_buf[359]*(20)+in_buf[360]*(2)+in_buf[361]*(0)+in_buf[362]*(-19)+in_buf[363]*(43)+in_buf[364]*(18)+in_buf[365]*(1)+in_buf[366]*(5)+in_buf[367]*(2)+in_buf[368]*(-27)+in_buf[369]*(0)+in_buf[370]*(-21)+in_buf[371]*(-30)+in_buf[372]*(-9)+in_buf[373]*(-15)+in_buf[374]*(-17)+in_buf[375]*(-10)+in_buf[376]*(0)+in_buf[377]*(16)+in_buf[378]*(28)+in_buf[379]*(22)+in_buf[380]*(10)+in_buf[381]*(-3)+in_buf[382]*(4)+in_buf[383]*(1)+in_buf[384]*(3)+in_buf[385]*(15)+in_buf[386]*(13)+in_buf[387]*(23)+in_buf[388]*(4)+in_buf[389]*(0)+in_buf[390]*(-8)+in_buf[391]*(2)+in_buf[392]*(3)+in_buf[393]*(-4)+in_buf[394]*(15)+in_buf[395]*(15)+in_buf[396]*(-31)+in_buf[397]*(-4)+in_buf[398]*(-10)+in_buf[399]*(-14)+in_buf[400]*(-34)+in_buf[401]*(-28)+in_buf[402]*(-26)+in_buf[403]*(-4)+in_buf[404]*(13)+in_buf[405]*(21)+in_buf[406]*(30)+in_buf[407]*(15)+in_buf[408]*(13)+in_buf[409]*(-17)+in_buf[410]*(-25)+in_buf[411]*(8)+in_buf[412]*(-2)+in_buf[413]*(-4)+in_buf[414]*(4)+in_buf[415]*(10)+in_buf[416]*(7)+in_buf[417]*(17)+in_buf[418]*(30)+in_buf[419]*(26)+in_buf[420]*(-2)+in_buf[421]*(-4)+in_buf[422]*(20)+in_buf[423]*(16)+in_buf[424]*(-36)+in_buf[425]*(-19)+in_buf[426]*(-22)+in_buf[427]*(-19)+in_buf[428]*(-27)+in_buf[429]*(-18)+in_buf[430]*(-4)+in_buf[431]*(24)+in_buf[432]*(31)+in_buf[433]*(36)+in_buf[434]*(28)+in_buf[435]*(8)+in_buf[436]*(-6)+in_buf[437]*(-27)+in_buf[438]*(-21)+in_buf[439]*(-8)+in_buf[440]*(-4)+in_buf[441]*(-6)+in_buf[442]*(-4)+in_buf[443]*(18)+in_buf[444]*(9)+in_buf[445]*(25)+in_buf[446]*(-14)+in_buf[447]*(28)+in_buf[448]*(-1)+in_buf[449]*(-5)+in_buf[450]*(8)+in_buf[451]*(-6)+in_buf[452]*(-25)+in_buf[453]*(-17)+in_buf[454]*(-25)+in_buf[455]*(-34)+in_buf[456]*(-16)+in_buf[457]*(8)+in_buf[458]*(29)+in_buf[459]*(51)+in_buf[460]*(52)+in_buf[461]*(34)+in_buf[462]*(13)+in_buf[463]*(-16)+in_buf[464]*(-9)+in_buf[465]*(-13)+in_buf[466]*(-1)+in_buf[467]*(-3)+in_buf[468]*(7)+in_buf[469]*(3)+in_buf[470]*(-10)+in_buf[471]*(-4)+in_buf[472]*(11)+in_buf[473]*(22)+in_buf[474]*(24)+in_buf[475]*(23)+in_buf[476]*(-2)+in_buf[477]*(-4)+in_buf[478]*(-3)+in_buf[479]*(-18)+in_buf[480]*(-30)+in_buf[481]*(-43)+in_buf[482]*(-26)+in_buf[483]*(-34)+in_buf[484]*(-19)+in_buf[485]*(17)+in_buf[486]*(42)+in_buf[487]*(45)+in_buf[488]*(44)+in_buf[489]*(18)+in_buf[490]*(-3)+in_buf[491]*(-34)+in_buf[492]*(-26)+in_buf[493]*(-29)+in_buf[494]*(-15)+in_buf[495]*(-6)+in_buf[496]*(9)+in_buf[497]*(-1)+in_buf[498]*(8)+in_buf[499]*(0)+in_buf[500]*(18)+in_buf[501]*(26)+in_buf[502]*(12)+in_buf[503]*(32)+in_buf[504]*(2)+in_buf[505]*(3)+in_buf[506]*(0)+in_buf[507]*(-20)+in_buf[508]*(-48)+in_buf[509]*(-53)+in_buf[510]*(-48)+in_buf[511]*(-19)+in_buf[512]*(-2)+in_buf[513]*(37)+in_buf[514]*(39)+in_buf[515]*(31)+in_buf[516]*(31)+in_buf[517]*(5)+in_buf[518]*(-21)+in_buf[519]*(-36)+in_buf[520]*(-30)+in_buf[521]*(-17)+in_buf[522]*(-18)+in_buf[523]*(-8)+in_buf[524]*(18)+in_buf[525]*(6)+in_buf[526]*(-1)+in_buf[527]*(9)+in_buf[528]*(9)+in_buf[529]*(51)+in_buf[530]*(29)+in_buf[531]*(37)+in_buf[532]*(22)+in_buf[533]*(-20)+in_buf[534]*(-18)+in_buf[535]*(4)+in_buf[536]*(-32)+in_buf[537]*(-48)+in_buf[538]*(-33)+in_buf[539]*(-16)+in_buf[540]*(-2)+in_buf[541]*(35)+in_buf[542]*(36)+in_buf[543]*(43)+in_buf[544]*(19)+in_buf[545]*(-1)+in_buf[546]*(-32)+in_buf[547]*(-35)+in_buf[548]*(-24)+in_buf[549]*(-17)+in_buf[550]*(-11)+in_buf[551]*(-10)+in_buf[552]*(8)+in_buf[553]*(-4)+in_buf[554]*(1)+in_buf[555]*(20)+in_buf[556]*(22)+in_buf[557]*(38)+in_buf[558]*(46)+in_buf[559]*(42)+in_buf[560]*(0)+in_buf[561]*(-24)+in_buf[562]*(-19)+in_buf[563]*(-12)+in_buf[564]*(-23)+in_buf[565]*(-26)+in_buf[566]*(-7)+in_buf[567]*(-8)+in_buf[568]*(-3)+in_buf[569]*(14)+in_buf[570]*(30)+in_buf[571]*(31)+in_buf[572]*(31)+in_buf[573]*(-10)+in_buf[574]*(-18)+in_buf[575]*(-18)+in_buf[576]*(-21)+in_buf[577]*(-11)+in_buf[578]*(-1)+in_buf[579]*(-6)+in_buf[580]*(1)+in_buf[581]*(-6)+in_buf[582]*(6)+in_buf[583]*(19)+in_buf[584]*(17)+in_buf[585]*(15)+in_buf[586]*(39)+in_buf[587]*(21)+in_buf[588]*(25)+in_buf[589]*(1)+in_buf[590]*(-2)+in_buf[591]*(-10)+in_buf[592]*(-17)+in_buf[593]*(7)+in_buf[594]*(14)+in_buf[595]*(0)+in_buf[596]*(-6)+in_buf[597]*(13)+in_buf[598]*(19)+in_buf[599]*(1)+in_buf[600]*(9)+in_buf[601]*(-7)+in_buf[602]*(-10)+in_buf[603]*(-14)+in_buf[604]*(-14)+in_buf[605]*(-12)+in_buf[606]*(-13)+in_buf[607]*(0)+in_buf[608]*(-1)+in_buf[609]*(3)+in_buf[610]*(11)+in_buf[611]*(32)+in_buf[612]*(-3)+in_buf[613]*(-8)+in_buf[614]*(26)+in_buf[615]*(-4)+in_buf[616]*(22)+in_buf[617]*(17)+in_buf[618]*(5)+in_buf[619]*(-21)+in_buf[620]*(8)+in_buf[621]*(44)+in_buf[622]*(10)+in_buf[623]*(11)+in_buf[624]*(6)+in_buf[625]*(5)+in_buf[626]*(7)+in_buf[627]*(-12)+in_buf[628]*(-8)+in_buf[629]*(-3)+in_buf[630]*(-7)+in_buf[631]*(3)+in_buf[632]*(2)+in_buf[633]*(-15)+in_buf[634]*(-12)+in_buf[635]*(-3)+in_buf[636]*(13)+in_buf[637]*(20)+in_buf[638]*(5)+in_buf[639]*(11)+in_buf[640]*(-15)+in_buf[641]*(-19)+in_buf[642]*(-11)+in_buf[643]*(-1)+in_buf[644]*(0)+in_buf[645]*(1)+in_buf[646]*(3)+in_buf[647]*(-37)+in_buf[648]*(-20)+in_buf[649]*(-6)+in_buf[650]*(-4)+in_buf[651]*(-7)+in_buf[652]*(-11)+in_buf[653]*(10)+in_buf[654]*(3)+in_buf[655]*(6)+in_buf[656]*(27)+in_buf[657]*(25)+in_buf[658]*(2)+in_buf[659]*(9)+in_buf[660]*(21)+in_buf[661]*(0)+in_buf[662]*(8)+in_buf[663]*(14)+in_buf[664]*(19)+in_buf[665]*(-3)+in_buf[666]*(-15)+in_buf[667]*(-13)+in_buf[668]*(-23)+in_buf[669]*(-16)+in_buf[670]*(0)+in_buf[671]*(2)+in_buf[672]*(2)+in_buf[673]*(3)+in_buf[674]*(-1)+in_buf[675]*(-37)+in_buf[676]*(-2)+in_buf[677]*(-2)+in_buf[678]*(-1)+in_buf[679]*(-24)+in_buf[680]*(-19)+in_buf[681]*(-2)+in_buf[682]*(14)+in_buf[683]*(25)+in_buf[684]*(24)+in_buf[685]*(0)+in_buf[686]*(7)+in_buf[687]*(2)+in_buf[688]*(-4)+in_buf[689]*(-30)+in_buf[690]*(-15)+in_buf[691]*(-10)+in_buf[692]*(-28)+in_buf[693]*(-41)+in_buf[694]*(-35)+in_buf[695]*(-19)+in_buf[696]*(11)+in_buf[697]*(35)+in_buf[698]*(21)+in_buf[699]*(4)+in_buf[700]*(-3)+in_buf[701]*(3)+in_buf[702]*(2)+in_buf[703]*(32)+in_buf[704]*(39)+in_buf[705]*(8)+in_buf[706]*(15)+in_buf[707]*(9)+in_buf[708]*(-13)+in_buf[709]*(0)+in_buf[710]*(2)+in_buf[711]*(0)+in_buf[712]*(-28)+in_buf[713]*(-19)+in_buf[714]*(0)+in_buf[715]*(-30)+in_buf[716]*(-46)+in_buf[717]*(-30)+in_buf[718]*(-49)+in_buf[719]*(-75)+in_buf[720]*(-60)+in_buf[721]*(-29)+in_buf[722]*(-38)+in_buf[723]*(-10)+in_buf[724]*(22)+in_buf[725]*(15)+in_buf[726]*(22)+in_buf[727]*(2)+in_buf[728]*(0)+in_buf[729]*(-3)+in_buf[730]*(3)+in_buf[731]*(-13)+in_buf[732]*(-19)+in_buf[733]*(35)+in_buf[734]*(48)+in_buf[735]*(40)+in_buf[736]*(-8)+in_buf[737]*(-39)+in_buf[738]*(-32)+in_buf[739]*(-18)+in_buf[740]*(-25)+in_buf[741]*(-43)+in_buf[742]*(-53)+in_buf[743]*(-55)+in_buf[744]*(-46)+in_buf[745]*(-26)+in_buf[746]*(-45)+in_buf[747]*(-51)+in_buf[748]*(-16)+in_buf[749]*(9)+in_buf[750]*(18)+in_buf[751]*(2)+in_buf[752]*(-2)+in_buf[753]*(4)+in_buf[754]*(-2)+in_buf[755]*(-2)+in_buf[756]*(1)+in_buf[757]*(1)+in_buf[758]*(0)+in_buf[759]*(2)+in_buf[760]*(21)+in_buf[761]*(19)+in_buf[762]*(24)+in_buf[763]*(1)+in_buf[764]*(-2)+in_buf[765]*(2)+in_buf[766]*(14)+in_buf[767]*(11)+in_buf[768]*(-14)+in_buf[769]*(-9)+in_buf[770]*(-3)+in_buf[771]*(8)+in_buf[772]*(4)+in_buf[773]*(-25)+in_buf[774]*(-23)+in_buf[775]*(-18)+in_buf[776]*(12)+in_buf[777]*(11)+in_buf[778]*(18)+in_buf[779]*(3)+in_buf[780]*(1)+in_buf[781]*(1)+in_buf[782]*(3)+in_buf[783]*(1);
assign in_buf_weight045=in_buf[0]*(3)+in_buf[1]*(0)+in_buf[2]*(-2)+in_buf[3]*(-2)+in_buf[4]*(0)+in_buf[5]*(-1)+in_buf[6]*(3)+in_buf[7]*(-2)+in_buf[8]*(4)+in_buf[9]*(-2)+in_buf[10]*(0)+in_buf[11]*(0)+in_buf[12]*(-5)+in_buf[13]*(-17)+in_buf[14]*(-15)+in_buf[15]*(-7)+in_buf[16]*(3)+in_buf[17]*(-3)+in_buf[18]*(3)+in_buf[19]*(-2)+in_buf[20]*(2)+in_buf[21]*(-1)+in_buf[22]*(1)+in_buf[23]*(0)+in_buf[24]*(-3)+in_buf[25]*(3)+in_buf[26]*(-1)+in_buf[27]*(-1)+in_buf[28]*(4)+in_buf[29]*(2)+in_buf[30]*(0)+in_buf[31]*(-4)+in_buf[32]*(-7)+in_buf[33]*(-1)+in_buf[34]*(0)+in_buf[35]*(0)+in_buf[36]*(-9)+in_buf[37]*(-6)+in_buf[38]*(11)+in_buf[39]*(-2)+in_buf[40]*(-16)+in_buf[41]*(-12)+in_buf[42]*(14)+in_buf[43]*(-32)+in_buf[44]*(-15)+in_buf[45]*(-23)+in_buf[46]*(-17)+in_buf[47]*(-14)+in_buf[48]*(-22)+in_buf[49]*(-26)+in_buf[50]*(-15)+in_buf[51]*(-4)+in_buf[52]*(-3)+in_buf[53]*(2)+in_buf[54]*(-1)+in_buf[55]*(-2)+in_buf[56]*(1)+in_buf[57]*(-2)+in_buf[58]*(-15)+in_buf[59]*(-29)+in_buf[60]*(-32)+in_buf[61]*(9)+in_buf[62]*(-1)+in_buf[63]*(-5)+in_buf[64]*(20)+in_buf[65]*(35)+in_buf[66]*(33)+in_buf[67]*(4)+in_buf[68]*(2)+in_buf[69]*(12)+in_buf[70]*(22)+in_buf[71]*(15)+in_buf[72]*(5)+in_buf[73]*(5)+in_buf[74]*(-10)+in_buf[75]*(-9)+in_buf[76]*(9)+in_buf[77]*(20)+in_buf[78]*(11)+in_buf[79]*(-4)+in_buf[80]*(13)+in_buf[81]*(5)+in_buf[82]*(-4)+in_buf[83]*(4)+in_buf[84]*(4)+in_buf[85]*(3)+in_buf[86]*(-12)+in_buf[87]*(-30)+in_buf[88]*(-35)+in_buf[89]*(0)+in_buf[90]*(0)+in_buf[91]*(-8)+in_buf[92]*(-13)+in_buf[93]*(17)+in_buf[94]*(5)+in_buf[95]*(14)+in_buf[96]*(0)+in_buf[97]*(5)+in_buf[98]*(0)+in_buf[99]*(10)+in_buf[100]*(8)+in_buf[101]*(-2)+in_buf[102]*(-6)+in_buf[103]*(-1)+in_buf[104]*(-35)+in_buf[105]*(-21)+in_buf[106]*(-5)+in_buf[107]*(-6)+in_buf[108]*(-4)+in_buf[109]*(-21)+in_buf[110]*(-1)+in_buf[111]*(0)+in_buf[112]*(0)+in_buf[113]*(-5)+in_buf[114]*(-20)+in_buf[115]*(-19)+in_buf[116]*(-9)+in_buf[117]*(-27)+in_buf[118]*(-13)+in_buf[119]*(-15)+in_buf[120]*(-4)+in_buf[121]*(3)+in_buf[122]*(13)+in_buf[123]*(2)+in_buf[124]*(13)+in_buf[125]*(12)+in_buf[126]*(16)+in_buf[127]*(-6)+in_buf[128]*(-4)+in_buf[129]*(-11)+in_buf[130]*(3)+in_buf[131]*(2)+in_buf[132]*(-3)+in_buf[133]*(-7)+in_buf[134]*(-6)+in_buf[135]*(-1)+in_buf[136]*(12)+in_buf[137]*(6)+in_buf[138]*(-36)+in_buf[139]*(16)+in_buf[140]*(-3)+in_buf[141]*(3)+in_buf[142]*(-30)+in_buf[143]*(20)+in_buf[144]*(21)+in_buf[145]*(-23)+in_buf[146]*(-26)+in_buf[147]*(-22)+in_buf[148]*(-21)+in_buf[149]*(-20)+in_buf[150]*(-5)+in_buf[151]*(0)+in_buf[152]*(19)+in_buf[153]*(11)+in_buf[154]*(8)+in_buf[155]*(-8)+in_buf[156]*(0)+in_buf[157]*(3)+in_buf[158]*(3)+in_buf[159]*(14)+in_buf[160]*(24)+in_buf[161]*(25)+in_buf[162]*(4)+in_buf[163]*(16)+in_buf[164]*(19)+in_buf[165]*(6)+in_buf[166]*(5)+in_buf[167]*(24)+in_buf[168]*(-3)+in_buf[169]*(1)+in_buf[170]*(14)+in_buf[171]*(14)+in_buf[172]*(27)+in_buf[173]*(-15)+in_buf[174]*(-27)+in_buf[175]*(-23)+in_buf[176]*(-37)+in_buf[177]*(-26)+in_buf[178]*(-24)+in_buf[179]*(0)+in_buf[180]*(23)+in_buf[181]*(13)+in_buf[182]*(-7)+in_buf[183]*(-21)+in_buf[184]*(-20)+in_buf[185]*(-23)+in_buf[186]*(-22)+in_buf[187]*(6)+in_buf[188]*(8)+in_buf[189]*(3)+in_buf[190]*(0)+in_buf[191]*(15)+in_buf[192]*(-3)+in_buf[193]*(2)+in_buf[194]*(8)+in_buf[195]*(19)+in_buf[196]*(-7)+in_buf[197]*(-9)+in_buf[198]*(22)+in_buf[199]*(4)+in_buf[200]*(19)+in_buf[201]*(-2)+in_buf[202]*(-6)+in_buf[203]*(-10)+in_buf[204]*(-15)+in_buf[205]*(-29)+in_buf[206]*(-25)+in_buf[207]*(12)+in_buf[208]*(20)+in_buf[209]*(7)+in_buf[210]*(-5)+in_buf[211]*(-34)+in_buf[212]*(-34)+in_buf[213]*(-13)+in_buf[214]*(-4)+in_buf[215]*(-3)+in_buf[216]*(-5)+in_buf[217]*(-7)+in_buf[218]*(3)+in_buf[219]*(-14)+in_buf[220]*(-9)+in_buf[221]*(-18)+in_buf[222]*(2)+in_buf[223]*(19)+in_buf[224]*(23)+in_buf[225]*(-26)+in_buf[226]*(16)+in_buf[227]*(6)+in_buf[228]*(6)+in_buf[229]*(-3)+in_buf[230]*(0)+in_buf[231]*(-9)+in_buf[232]*(-29)+in_buf[233]*(-16)+in_buf[234]*(-12)+in_buf[235]*(13)+in_buf[236]*(19)+in_buf[237]*(17)+in_buf[238]*(-9)+in_buf[239]*(-17)+in_buf[240]*(-26)+in_buf[241]*(-6)+in_buf[242]*(0)+in_buf[243]*(7)+in_buf[244]*(-13)+in_buf[245]*(-13)+in_buf[246]*(-17)+in_buf[247]*(-22)+in_buf[248]*(-28)+in_buf[249]*(-36)+in_buf[250]*(-9)+in_buf[251]*(-10)+in_buf[252]*(-15)+in_buf[253]*(-34)+in_buf[254]*(5)+in_buf[255]*(2)+in_buf[256]*(-6)+in_buf[257]*(5)+in_buf[258]*(-13)+in_buf[259]*(-17)+in_buf[260]*(-20)+in_buf[261]*(-21)+in_buf[262]*(-13)+in_buf[263]*(10)+in_buf[264]*(15)+in_buf[265]*(11)+in_buf[266]*(-11)+in_buf[267]*(-13)+in_buf[268]*(-13)+in_buf[269]*(-6)+in_buf[270]*(17)+in_buf[271]*(9)+in_buf[272]*(-2)+in_buf[273]*(-1)+in_buf[274]*(-14)+in_buf[275]*(-38)+in_buf[276]*(-30)+in_buf[277]*(-36)+in_buf[278]*(-10)+in_buf[279]*(-16)+in_buf[280]*(-13)+in_buf[281]*(-12)+in_buf[282]*(-1)+in_buf[283]*(16)+in_buf[284]*(9)+in_buf[285]*(18)+in_buf[286]*(-3)+in_buf[287]*(-15)+in_buf[288]*(-14)+in_buf[289]*(-22)+in_buf[290]*(-4)+in_buf[291]*(11)+in_buf[292]*(13)+in_buf[293]*(7)+in_buf[294]*(-8)+in_buf[295]*(-29)+in_buf[296]*(-17)+in_buf[297]*(18)+in_buf[298]*(15)+in_buf[299]*(0)+in_buf[300]*(-12)+in_buf[301]*(0)+in_buf[302]*(-16)+in_buf[303]*(-29)+in_buf[304]*(-23)+in_buf[305]*(-19)+in_buf[306]*(-5)+in_buf[307]*(-6)+in_buf[308]*(-17)+in_buf[309]*(5)+in_buf[310]*(-1)+in_buf[311]*(12)+in_buf[312]*(-1)+in_buf[313]*(-6)+in_buf[314]*(4)+in_buf[315]*(-5)+in_buf[316]*(-6)+in_buf[317]*(-23)+in_buf[318]*(1)+in_buf[319]*(-1)+in_buf[320]*(14)+in_buf[321]*(-8)+in_buf[322]*(-26)+in_buf[323]*(-36)+in_buf[324]*(-3)+in_buf[325]*(14)+in_buf[326]*(10)+in_buf[327]*(9)+in_buf[328]*(-28)+in_buf[329]*(-8)+in_buf[330]*(-1)+in_buf[331]*(-15)+in_buf[332]*(-7)+in_buf[333]*(4)+in_buf[334]*(-29)+in_buf[335]*(-18)+in_buf[336]*(-12)+in_buf[337]*(4)+in_buf[338]*(11)+in_buf[339]*(-4)+in_buf[340]*(-3)+in_buf[341]*(-13)+in_buf[342]*(-14)+in_buf[343]*(-15)+in_buf[344]*(-23)+in_buf[345]*(-17)+in_buf[346]*(-4)+in_buf[347]*(7)+in_buf[348]*(9)+in_buf[349]*(-15)+in_buf[350]*(-24)+in_buf[351]*(-30)+in_buf[352]*(-6)+in_buf[353]*(5)+in_buf[354]*(-4)+in_buf[355]*(-21)+in_buf[356]*(-17)+in_buf[357]*(-12)+in_buf[358]*(4)+in_buf[359]*(-13)+in_buf[360]*(28)+in_buf[361]*(23)+in_buf[362]*(-12)+in_buf[363]*(-22)+in_buf[364]*(-2)+in_buf[365]*(19)+in_buf[366]*(27)+in_buf[367]*(-21)+in_buf[368]*(-22)+in_buf[369]*(-12)+in_buf[370]*(-1)+in_buf[371]*(-18)+in_buf[372]*(-12)+in_buf[373]*(-10)+in_buf[374]*(2)+in_buf[375]*(11)+in_buf[376]*(5)+in_buf[377]*(-2)+in_buf[378]*(-22)+in_buf[379]*(-18)+in_buf[380]*(-11)+in_buf[381]*(2)+in_buf[382]*(-9)+in_buf[383]*(-16)+in_buf[384]*(-16)+in_buf[385]*(-3)+in_buf[386]*(0)+in_buf[387]*(0)+in_buf[388]*(25)+in_buf[389]*(35)+in_buf[390]*(16)+in_buf[391]*(19)+in_buf[392]*(1)+in_buf[393]*(12)+in_buf[394]*(27)+in_buf[395]*(-14)+in_buf[396]*(-3)+in_buf[397]*(-3)+in_buf[398]*(4)+in_buf[399]*(-1)+in_buf[400]*(-9)+in_buf[401]*(-1)+in_buf[402]*(-4)+in_buf[403]*(3)+in_buf[404]*(12)+in_buf[405]*(3)+in_buf[406]*(2)+in_buf[407]*(-6)+in_buf[408]*(6)+in_buf[409]*(-3)+in_buf[410]*(-13)+in_buf[411]*(-15)+in_buf[412]*(-20)+in_buf[413]*(-15)+in_buf[414]*(-2)+in_buf[415]*(-18)+in_buf[416]*(0)+in_buf[417]*(68)+in_buf[418]*(61)+in_buf[419]*(20)+in_buf[420]*(0)+in_buf[421]*(-2)+in_buf[422]*(28)+in_buf[423]*(27)+in_buf[424]*(18)+in_buf[425]*(19)+in_buf[426]*(11)+in_buf[427]*(2)+in_buf[428]*(4)+in_buf[429]*(9)+in_buf[430]*(4)+in_buf[431]*(5)+in_buf[432]*(17)+in_buf[433]*(21)+in_buf[434]*(5)+in_buf[435]*(12)+in_buf[436]*(16)+in_buf[437]*(10)+in_buf[438]*(-13)+in_buf[439]*(1)+in_buf[440]*(-16)+in_buf[441]*(-7)+in_buf[442]*(2)+in_buf[443]*(-11)+in_buf[444]*(-2)+in_buf[445]*(38)+in_buf[446]*(59)+in_buf[447]*(29)+in_buf[448]*(-5)+in_buf[449]*(-11)+in_buf[450]*(7)+in_buf[451]*(22)+in_buf[452]*(5)+in_buf[453]*(12)+in_buf[454]*(14)+in_buf[455]*(12)+in_buf[456]*(14)+in_buf[457]*(22)+in_buf[458]*(15)+in_buf[459]*(12)+in_buf[460]*(10)+in_buf[461]*(6)+in_buf[462]*(1)+in_buf[463]*(19)+in_buf[464]*(33)+in_buf[465]*(19)+in_buf[466]*(15)+in_buf[467]*(20)+in_buf[468]*(9)+in_buf[469]*(45)+in_buf[470]*(32)+in_buf[471]*(13)+in_buf[472]*(0)+in_buf[473]*(49)+in_buf[474]*(71)+in_buf[475]*(21)+in_buf[476]*(2)+in_buf[477]*(-5)+in_buf[478]*(25)+in_buf[479]*(4)+in_buf[480]*(14)+in_buf[481]*(11)+in_buf[482]*(16)+in_buf[483]*(15)+in_buf[484]*(21)+in_buf[485]*(16)+in_buf[486]*(4)+in_buf[487]*(0)+in_buf[488]*(-2)+in_buf[489]*(2)+in_buf[490]*(15)+in_buf[491]*(20)+in_buf[492]*(23)+in_buf[493]*(25)+in_buf[494]*(26)+in_buf[495]*(15)+in_buf[496]*(22)+in_buf[497]*(44)+in_buf[498]*(21)+in_buf[499]*(17)+in_buf[500]*(15)+in_buf[501]*(31)+in_buf[502]*(46)+in_buf[503]*(7)+in_buf[504]*(-31)+in_buf[505]*(-11)+in_buf[506]*(16)+in_buf[507]*(15)+in_buf[508]*(18)+in_buf[509]*(13)+in_buf[510]*(10)+in_buf[511]*(20)+in_buf[512]*(14)+in_buf[513]*(11)+in_buf[514]*(-1)+in_buf[515]*(-14)+in_buf[516]*(6)+in_buf[517]*(16)+in_buf[518]*(25)+in_buf[519]*(12)+in_buf[520]*(24)+in_buf[521]*(13)+in_buf[522]*(6)+in_buf[523]*(11)+in_buf[524]*(18)+in_buf[525]*(28)+in_buf[526]*(13)+in_buf[527]*(26)+in_buf[528]*(30)+in_buf[529]*(24)+in_buf[530]*(22)+in_buf[531]*(37)+in_buf[532]*(-3)+in_buf[533]*(-32)+in_buf[534]*(-7)+in_buf[535]*(24)+in_buf[536]*(17)+in_buf[537]*(12)+in_buf[538]*(1)+in_buf[539]*(10)+in_buf[540]*(7)+in_buf[541]*(14)+in_buf[542]*(14)+in_buf[543]*(0)+in_buf[544]*(-2)+in_buf[545]*(10)+in_buf[546]*(16)+in_buf[547]*(15)+in_buf[548]*(20)+in_buf[549]*(26)+in_buf[550]*(11)+in_buf[551]*(12)+in_buf[552]*(23)+in_buf[553]*(22)+in_buf[554]*(21)+in_buf[555]*(37)+in_buf[556]*(20)+in_buf[557]*(26)+in_buf[558]*(56)+in_buf[559]*(19)+in_buf[560]*(0)+in_buf[561]*(-2)+in_buf[562]*(6)+in_buf[563]*(29)+in_buf[564]*(4)+in_buf[565]*(-2)+in_buf[566]*(6)+in_buf[567]*(22)+in_buf[568]*(7)+in_buf[569]*(8)+in_buf[570]*(-2)+in_buf[571]*(-5)+in_buf[572]*(6)+in_buf[573]*(1)+in_buf[574]*(4)+in_buf[575]*(7)+in_buf[576]*(11)+in_buf[577]*(14)+in_buf[578]*(11)+in_buf[579]*(13)+in_buf[580]*(16)+in_buf[581]*(12)+in_buf[582]*(16)+in_buf[583]*(29)+in_buf[584]*(6)+in_buf[585]*(2)+in_buf[586]*(40)+in_buf[587]*(-6)+in_buf[588]*(0)+in_buf[589]*(7)+in_buf[590]*(-4)+in_buf[591]*(24)+in_buf[592]*(9)+in_buf[593]*(8)+in_buf[594]*(-3)+in_buf[595]*(5)+in_buf[596]*(9)+in_buf[597]*(9)+in_buf[598]*(-3)+in_buf[599]*(-14)+in_buf[600]*(-3)+in_buf[601]*(2)+in_buf[602]*(-6)+in_buf[603]*(-3)+in_buf[604]*(4)+in_buf[605]*(6)+in_buf[606]*(7)+in_buf[607]*(10)+in_buf[608]*(13)+in_buf[609]*(6)+in_buf[610]*(42)+in_buf[611]*(51)+in_buf[612]*(21)+in_buf[613]*(9)+in_buf[614]*(3)+in_buf[615]*(-1)+in_buf[616]*(-3)+in_buf[617]*(-1)+in_buf[618]*(5)+in_buf[619]*(5)+in_buf[620]*(15)+in_buf[621]*(23)+in_buf[622]*(-11)+in_buf[623]*(-13)+in_buf[624]*(-3)+in_buf[625]*(0)+in_buf[626]*(4)+in_buf[627]*(-4)+in_buf[628]*(-8)+in_buf[629]*(-9)+in_buf[630]*(-23)+in_buf[631]*(-14)+in_buf[632]*(-14)+in_buf[633]*(-11)+in_buf[634]*(-12)+in_buf[635]*(5)+in_buf[636]*(9)+in_buf[637]*(16)+in_buf[638]*(30)+in_buf[639]*(35)+in_buf[640]*(20)+in_buf[641]*(-11)+in_buf[642]*(-18)+in_buf[643]*(0)+in_buf[644]*(1)+in_buf[645]*(0)+in_buf[646]*(11)+in_buf[647]*(30)+in_buf[648]*(9)+in_buf[649]*(6)+in_buf[650]*(-3)+in_buf[651]*(-12)+in_buf[652]*(-2)+in_buf[653]*(-9)+in_buf[654]*(-10)+in_buf[655]*(2)+in_buf[656]*(5)+in_buf[657]*(-4)+in_buf[658]*(-11)+in_buf[659]*(0)+in_buf[660]*(0)+in_buf[661]*(-23)+in_buf[662]*(-3)+in_buf[663]*(-5)+in_buf[664]*(3)+in_buf[665]*(28)+in_buf[666]*(18)+in_buf[667]*(22)+in_buf[668]*(0)+in_buf[669]*(-9)+in_buf[670]*(-12)+in_buf[671]*(2)+in_buf[672]*(-3)+in_buf[673]*(0)+in_buf[674]*(2)+in_buf[675]*(-2)+in_buf[676]*(0)+in_buf[677]*(1)+in_buf[678]*(-18)+in_buf[679]*(-16)+in_buf[680]*(-19)+in_buf[681]*(-17)+in_buf[682]*(-17)+in_buf[683]*(-1)+in_buf[684]*(-23)+in_buf[685]*(-8)+in_buf[686]*(3)+in_buf[687]*(0)+in_buf[688]*(13)+in_buf[689]*(-14)+in_buf[690]*(-15)+in_buf[691]*(-26)+in_buf[692]*(-11)+in_buf[693]*(5)+in_buf[694]*(4)+in_buf[695]*(7)+in_buf[696]*(26)+in_buf[697]*(13)+in_buf[698]*(8)+in_buf[699]*(4)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(-1)+in_buf[703]*(-11)+in_buf[704]*(-13)+in_buf[705]*(-25)+in_buf[706]*(-25)+in_buf[707]*(-19)+in_buf[708]*(-30)+in_buf[709]*(-64)+in_buf[710]*(-36)+in_buf[711]*(-13)+in_buf[712]*(-58)+in_buf[713]*(-35)+in_buf[714]*(-37)+in_buf[715]*(-25)+in_buf[716]*(-9)+in_buf[717]*(-26)+in_buf[718]*(-28)+in_buf[719]*(-50)+in_buf[720]*(-48)+in_buf[721]*(-60)+in_buf[722]*(-35)+in_buf[723]*(-5)+in_buf[724]*(-12)+in_buf[725]*(-1)+in_buf[726]*(16)+in_buf[727]*(2)+in_buf[728]*(4)+in_buf[729]*(1)+in_buf[730]*(-1)+in_buf[731]*(-1)+in_buf[732]*(1)+in_buf[733]*(-6)+in_buf[734]*(-15)+in_buf[735]*(-28)+in_buf[736]*(-38)+in_buf[737]*(-55)+in_buf[738]*(-42)+in_buf[739]*(-53)+in_buf[740]*(-51)+in_buf[741]*(-51)+in_buf[742]*(-82)+in_buf[743]*(-69)+in_buf[744]*(-41)+in_buf[745]*(-34)+in_buf[746]*(-42)+in_buf[747]*(-44)+in_buf[748]*(-42)+in_buf[749]*(-35)+in_buf[750]*(-17)+in_buf[751]*(13)+in_buf[752]*(-12)+in_buf[753]*(2)+in_buf[754]*(1)+in_buf[755]*(1)+in_buf[756]*(-2)+in_buf[757]*(-2)+in_buf[758]*(-3)+in_buf[759]*(4)+in_buf[760]*(-3)+in_buf[761]*(0)+in_buf[762]*(-6)+in_buf[763]*(-6)+in_buf[764]*(-13)+in_buf[765]*(-4)+in_buf[766]*(-31)+in_buf[767]*(-22)+in_buf[768]*(-16)+in_buf[769]*(-22)+in_buf[770]*(-40)+in_buf[771]*(-7)+in_buf[772]*(-5)+in_buf[773]*(-33)+in_buf[774]*(-41)+in_buf[775]*(-15)+in_buf[776]*(0)+in_buf[777]*(-15)+in_buf[778]*(-22)+in_buf[779]*(-16)+in_buf[780]*(4)+in_buf[781]*(4)+in_buf[782]*(-1)+in_buf[783]*(3);
assign in_buf_weight046=in_buf[0]*(2)+in_buf[1]*(-2)+in_buf[2]*(2)+in_buf[3]*(4)+in_buf[4]*(1)+in_buf[5]*(3)+in_buf[6]*(2)+in_buf[7]*(2)+in_buf[8]*(0)+in_buf[9]*(-1)+in_buf[10]*(2)+in_buf[11]*(3)+in_buf[12]*(0)+in_buf[13]*(-2)+in_buf[14]*(0)+in_buf[15]*(0)+in_buf[16]*(0)+in_buf[17]*(3)+in_buf[18]*(0)+in_buf[19]*(3)+in_buf[20]*(2)+in_buf[21]*(3)+in_buf[22]*(3)+in_buf[23]*(1)+in_buf[24]*(1)+in_buf[25]*(2)+in_buf[26]*(-2)+in_buf[27]*(2)+in_buf[28]*(1)+in_buf[29]*(-1)+in_buf[30]*(-3)+in_buf[31]*(-2)+in_buf[32]*(-4)+in_buf[33]*(0)+in_buf[34]*(-10)+in_buf[35]*(-10)+in_buf[36]*(-8)+in_buf[37]*(-6)+in_buf[38]*(-13)+in_buf[39]*(-20)+in_buf[40]*(-12)+in_buf[41]*(-27)+in_buf[42]*(-20)+in_buf[43]*(-2)+in_buf[44]*(10)+in_buf[45]*(-2)+in_buf[46]*(-6)+in_buf[47]*(-11)+in_buf[48]*(-20)+in_buf[49]*(-8)+in_buf[50]*(0)+in_buf[51]*(-5)+in_buf[52]*(4)+in_buf[53]*(1)+in_buf[54]*(0)+in_buf[55]*(4)+in_buf[56]*(2)+in_buf[57]*(0)+in_buf[58]*(1)+in_buf[59]*(1)+in_buf[60]*(-6)+in_buf[61]*(-5)+in_buf[62]*(-7)+in_buf[63]*(-8)+in_buf[64]*(22)+in_buf[65]*(18)+in_buf[66]*(10)+in_buf[67]*(10)+in_buf[68]*(6)+in_buf[69]*(-24)+in_buf[70]*(-9)+in_buf[71]*(3)+in_buf[72]*(7)+in_buf[73]*(16)+in_buf[74]*(23)+in_buf[75]*(10)+in_buf[76]*(-11)+in_buf[77]*(-7)+in_buf[78]*(0)+in_buf[79]*(19)+in_buf[80]*(15)+in_buf[81]*(3)+in_buf[82]*(-1)+in_buf[83]*(-1)+in_buf[84]*(3)+in_buf[85]*(2)+in_buf[86]*(-14)+in_buf[87]*(-3)+in_buf[88]*(-2)+in_buf[89]*(1)+in_buf[90]*(12)+in_buf[91]*(0)+in_buf[92]*(-12)+in_buf[93]*(3)+in_buf[94]*(-3)+in_buf[95]*(-10)+in_buf[96]*(-35)+in_buf[97]*(-44)+in_buf[98]*(-52)+in_buf[99]*(-28)+in_buf[100]*(-5)+in_buf[101]*(-22)+in_buf[102]*(-35)+in_buf[103]*(-9)+in_buf[104]*(-39)+in_buf[105]*(-15)+in_buf[106]*(-15)+in_buf[107]*(10)+in_buf[108]*(20)+in_buf[109]*(12)+in_buf[110]*(-5)+in_buf[111]*(-2)+in_buf[112]*(3)+in_buf[113]*(-1)+in_buf[114]*(-7)+in_buf[115]*(-17)+in_buf[116]*(11)+in_buf[117]*(5)+in_buf[118]*(0)+in_buf[119]*(6)+in_buf[120]*(12)+in_buf[121]*(16)+in_buf[122]*(3)+in_buf[123]*(-1)+in_buf[124]*(-16)+in_buf[125]*(-38)+in_buf[126]*(-45)+in_buf[127]*(-45)+in_buf[128]*(-28)+in_buf[129]*(-7)+in_buf[130]*(-21)+in_buf[131]*(-13)+in_buf[132]*(-5)+in_buf[133]*(4)+in_buf[134]*(-4)+in_buf[135]*(-22)+in_buf[136]*(-7)+in_buf[137]*(33)+in_buf[138]*(37)+in_buf[139]*(11)+in_buf[140]*(-1)+in_buf[141]*(-1)+in_buf[142]*(-8)+in_buf[143]*(12)+in_buf[144]*(32)+in_buf[145]*(-2)+in_buf[146]*(-10)+in_buf[147]*(13)+in_buf[148]*(31)+in_buf[149]*(13)+in_buf[150]*(11)+in_buf[151]*(16)+in_buf[152]*(15)+in_buf[153]*(4)+in_buf[154]*(-15)+in_buf[155]*(-13)+in_buf[156]*(-12)+in_buf[157]*(-10)+in_buf[158]*(-14)+in_buf[159]*(-8)+in_buf[160]*(0)+in_buf[161]*(7)+in_buf[162]*(1)+in_buf[163]*(5)+in_buf[164]*(7)+in_buf[165]*(33)+in_buf[166]*(18)+in_buf[167]*(-3)+in_buf[168]*(0)+in_buf[169]*(0)+in_buf[170]*(4)+in_buf[171]*(28)+in_buf[172]*(25)+in_buf[173]*(-3)+in_buf[174]*(8)+in_buf[175]*(13)+in_buf[176]*(16)+in_buf[177]*(20)+in_buf[178]*(11)+in_buf[179]*(-3)+in_buf[180]*(14)+in_buf[181]*(4)+in_buf[182]*(0)+in_buf[183]*(-4)+in_buf[184]*(11)+in_buf[185]*(11)+in_buf[186]*(-2)+in_buf[187]*(0)+in_buf[188]*(12)+in_buf[189]*(29)+in_buf[190]*(6)+in_buf[191]*(27)+in_buf[192]*(-1)+in_buf[193]*(-6)+in_buf[194]*(-8)+in_buf[195]*(-4)+in_buf[196]*(1)+in_buf[197]*(0)+in_buf[198]*(31)+in_buf[199]*(29)+in_buf[200]*(16)+in_buf[201]*(-13)+in_buf[202]*(2)+in_buf[203]*(8)+in_buf[204]*(3)+in_buf[205]*(2)+in_buf[206]*(-4)+in_buf[207]*(-2)+in_buf[208]*(-8)+in_buf[209]*(2)+in_buf[210]*(-10)+in_buf[211]*(-6)+in_buf[212]*(-6)+in_buf[213]*(2)+in_buf[214]*(6)+in_buf[215]*(-7)+in_buf[216]*(-2)+in_buf[217]*(22)+in_buf[218]*(19)+in_buf[219]*(12)+in_buf[220]*(1)+in_buf[221]*(0)+in_buf[222]*(-4)+in_buf[223]*(-22)+in_buf[224]*(3)+in_buf[225]*(20)+in_buf[226]*(20)+in_buf[227]*(12)+in_buf[228]*(22)+in_buf[229]*(12)+in_buf[230]*(10)+in_buf[231]*(9)+in_buf[232]*(18)+in_buf[233]*(-3)+in_buf[234]*(-1)+in_buf[235]*(-7)+in_buf[236]*(9)+in_buf[237]*(17)+in_buf[238]*(7)+in_buf[239]*(0)+in_buf[240]*(-5)+in_buf[241]*(-11)+in_buf[242]*(3)+in_buf[243]*(0)+in_buf[244]*(-4)+in_buf[245]*(-1)+in_buf[246]*(-4)+in_buf[247]*(27)+in_buf[248]*(3)+in_buf[249]*(19)+in_buf[250]*(29)+in_buf[251]*(0)+in_buf[252]*(6)+in_buf[253]*(30)+in_buf[254]*(16)+in_buf[255]*(27)+in_buf[256]*(8)+in_buf[257]*(36)+in_buf[258]*(5)+in_buf[259]*(-6)+in_buf[260]*(0)+in_buf[261]*(-3)+in_buf[262]*(3)+in_buf[263]*(2)+in_buf[264]*(29)+in_buf[265]*(21)+in_buf[266]*(-1)+in_buf[267]*(-7)+in_buf[268]*(-12)+in_buf[269]*(3)+in_buf[270]*(9)+in_buf[271]*(3)+in_buf[272]*(-1)+in_buf[273]*(-7)+in_buf[274]*(-7)+in_buf[275]*(5)+in_buf[276]*(-5)+in_buf[277]*(47)+in_buf[278]*(41)+in_buf[279]*(26)+in_buf[280]*(16)+in_buf[281]*(12)+in_buf[282]*(21)+in_buf[283]*(10)+in_buf[284]*(5)+in_buf[285]*(37)+in_buf[286]*(27)+in_buf[287]*(-4)+in_buf[288]*(-3)+in_buf[289]*(5)+in_buf[290]*(19)+in_buf[291]*(26)+in_buf[292]*(13)+in_buf[293]*(6)+in_buf[294]*(-25)+in_buf[295]*(-19)+in_buf[296]*(4)+in_buf[297]*(9)+in_buf[298]*(6)+in_buf[299]*(4)+in_buf[300]*(-5)+in_buf[301]*(-7)+in_buf[302]*(-9)+in_buf[303]*(4)+in_buf[304]*(33)+in_buf[305]*(14)+in_buf[306]*(-25)+in_buf[307]*(27)+in_buf[308]*(9)+in_buf[309]*(35)+in_buf[310]*(-2)+in_buf[311]*(9)+in_buf[312]*(4)+in_buf[313]*(21)+in_buf[314]*(29)+in_buf[315]*(23)+in_buf[316]*(16)+in_buf[317]*(20)+in_buf[318]*(20)+in_buf[319]*(28)+in_buf[320]*(4)+in_buf[321]*(-22)+in_buf[322]*(-42)+in_buf[323]*(-14)+in_buf[324]*(15)+in_buf[325]*(11)+in_buf[326]*(0)+in_buf[327]*(5)+in_buf[328]*(9)+in_buf[329]*(-3)+in_buf[330]*(-12)+in_buf[331]*(10)+in_buf[332]*(32)+in_buf[333]*(3)+in_buf[334]*(-36)+in_buf[335]*(-24)+in_buf[336]*(8)+in_buf[337]*(10)+in_buf[338]*(-1)+in_buf[339]*(-8)+in_buf[340]*(16)+in_buf[341]*(15)+in_buf[342]*(8)+in_buf[343]*(10)+in_buf[344]*(10)+in_buf[345]*(12)+in_buf[346]*(2)+in_buf[347]*(-7)+in_buf[348]*(-18)+in_buf[349]*(-46)+in_buf[350]*(-36)+in_buf[351]*(-1)+in_buf[352]*(18)+in_buf[353]*(11)+in_buf[354]*(-3)+in_buf[355]*(1)+in_buf[356]*(-8)+in_buf[357]*(-10)+in_buf[358]*(-4)+in_buf[359]*(-22)+in_buf[360]*(1)+in_buf[361]*(0)+in_buf[362]*(-23)+in_buf[363]*(-14)+in_buf[364]*(-15)+in_buf[365]*(28)+in_buf[366]*(47)+in_buf[367]*(-4)+in_buf[368]*(-6)+in_buf[369]*(0)+in_buf[370]*(8)+in_buf[371]*(4)+in_buf[372]*(-2)+in_buf[373]*(2)+in_buf[374]*(-11)+in_buf[375]*(-26)+in_buf[376]*(-53)+in_buf[377]*(-33)+in_buf[378]*(-8)+in_buf[379]*(0)+in_buf[380]*(12)+in_buf[381]*(15)+in_buf[382]*(7)+in_buf[383]*(-4)+in_buf[384]*(-17)+in_buf[385]*(4)+in_buf[386]*(7)+in_buf[387]*(-4)+in_buf[388]*(-16)+in_buf[389]*(2)+in_buf[390]*(24)+in_buf[391]*(5)+in_buf[392]*(-15)+in_buf[393]*(23)+in_buf[394]*(32)+in_buf[395]*(1)+in_buf[396]*(-15)+in_buf[397]*(1)+in_buf[398]*(9)+in_buf[399]*(-9)+in_buf[400]*(-22)+in_buf[401]*(-24)+in_buf[402]*(-30)+in_buf[403]*(-46)+in_buf[404]*(-28)+in_buf[405]*(-10)+in_buf[406]*(-1)+in_buf[407]*(14)+in_buf[408]*(9)+in_buf[409]*(8)+in_buf[410]*(-1)+in_buf[411]*(18)+in_buf[412]*(-5)+in_buf[413]*(-11)+in_buf[414]*(-12)+in_buf[415]*(0)+in_buf[416]*(-13)+in_buf[417]*(7)+in_buf[418]*(30)+in_buf[419]*(13)+in_buf[420]*(-9)+in_buf[421]*(2)+in_buf[422]*(9)+in_buf[423]*(-18)+in_buf[424]*(-11)+in_buf[425]*(-13)+in_buf[426]*(-16)+in_buf[427]*(-32)+in_buf[428]*(-44)+in_buf[429]*(-44)+in_buf[430]*(-54)+in_buf[431]*(-35)+in_buf[432]*(-11)+in_buf[433]*(13)+in_buf[434]*(27)+in_buf[435]*(22)+in_buf[436]*(2)+in_buf[437]*(3)+in_buf[438]*(3)+in_buf[439]*(16)+in_buf[440]*(7)+in_buf[441]*(-15)+in_buf[442]*(-17)+in_buf[443]*(-15)+in_buf[444]*(-18)+in_buf[445]*(-14)+in_buf[446]*(0)+in_buf[447]*(12)+in_buf[448]*(10)+in_buf[449]*(-8)+in_buf[450]*(-3)+in_buf[451]*(-28)+in_buf[452]*(-15)+in_buf[453]*(-31)+in_buf[454]*(-40)+in_buf[455]*(-75)+in_buf[456]*(-93)+in_buf[457]*(-89)+in_buf[458]*(-42)+in_buf[459]*(1)+in_buf[460]*(21)+in_buf[461]*(15)+in_buf[462]*(19)+in_buf[463]*(10)+in_buf[464]*(14)+in_buf[465]*(8)+in_buf[466]*(8)+in_buf[467]*(10)+in_buf[468]*(0)+in_buf[469]*(2)+in_buf[470]*(0)+in_buf[471]*(2)+in_buf[472]*(-8)+in_buf[473]*(-2)+in_buf[474]*(0)+in_buf[475]*(10)+in_buf[476]*(-3)+in_buf[477]*(-4)+in_buf[478]*(-2)+in_buf[479]*(-20)+in_buf[480]*(-37)+in_buf[481]*(-24)+in_buf[482]*(-61)+in_buf[483]*(-83)+in_buf[484]*(-75)+in_buf[485]*(-52)+in_buf[486]*(-22)+in_buf[487]*(30)+in_buf[488]*(33)+in_buf[489]*(19)+in_buf[490]*(16)+in_buf[491]*(10)+in_buf[492]*(4)+in_buf[493]*(4)+in_buf[494]*(13)+in_buf[495]*(13)+in_buf[496]*(-2)+in_buf[497]*(-12)+in_buf[498]*(-3)+in_buf[499]*(4)+in_buf[500]*(26)+in_buf[501]*(28)+in_buf[502]*(1)+in_buf[503]*(21)+in_buf[504]*(13)+in_buf[505]*(-8)+in_buf[506]*(0)+in_buf[507]*(-17)+in_buf[508]*(-22)+in_buf[509]*(-35)+in_buf[510]*(-48)+in_buf[511]*(-50)+in_buf[512]*(-36)+in_buf[513]*(-16)+in_buf[514]*(20)+in_buf[515]*(37)+in_buf[516]*(28)+in_buf[517]*(22)+in_buf[518]*(5)+in_buf[519]*(10)+in_buf[520]*(-5)+in_buf[521]*(2)+in_buf[522]*(1)+in_buf[523]*(-12)+in_buf[524]*(-18)+in_buf[525]*(-30)+in_buf[526]*(-7)+in_buf[527]*(-2)+in_buf[528]*(5)+in_buf[529]*(23)+in_buf[530]*(-6)+in_buf[531]*(1)+in_buf[532]*(-18)+in_buf[533]*(16)+in_buf[534]*(-8)+in_buf[535]*(-26)+in_buf[536]*(-27)+in_buf[537]*(-44)+in_buf[538]*(-55)+in_buf[539]*(-29)+in_buf[540]*(-6)+in_buf[541]*(18)+in_buf[542]*(39)+in_buf[543]*(29)+in_buf[544]*(19)+in_buf[545]*(8)+in_buf[546]*(4)+in_buf[547]*(5)+in_buf[548]*(5)+in_buf[549]*(5)+in_buf[550]*(-7)+in_buf[551]*(-7)+in_buf[552]*(-4)+in_buf[553]*(-18)+in_buf[554]*(-6)+in_buf[555]*(0)+in_buf[556]*(-3)+in_buf[557]*(22)+in_buf[558]*(36)+in_buf[559]*(-21)+in_buf[560]*(-2)+in_buf[561]*(-6)+in_buf[562]*(-17)+in_buf[563]*(-25)+in_buf[564]*(-46)+in_buf[565]*(-48)+in_buf[566]*(-32)+in_buf[567]*(-15)+in_buf[568]*(8)+in_buf[569]*(16)+in_buf[570]*(29)+in_buf[571]*(25)+in_buf[572]*(20)+in_buf[573]*(3)+in_buf[574]*(-8)+in_buf[575]*(8)+in_buf[576]*(11)+in_buf[577]*(-3)+in_buf[578]*(-20)+in_buf[579]*(-8)+in_buf[580]*(7)+in_buf[581]*(0)+in_buf[582]*(-8)+in_buf[583]*(-14)+in_buf[584]*(17)+in_buf[585]*(42)+in_buf[586]*(34)+in_buf[587]*(-16)+in_buf[588]*(-22)+in_buf[589]*(0)+in_buf[590]*(-13)+in_buf[591]*(-35)+in_buf[592]*(-57)+in_buf[593]*(-41)+in_buf[594]*(-30)+in_buf[595]*(-23)+in_buf[596]*(-13)+in_buf[597]*(15)+in_buf[598]*(8)+in_buf[599]*(4)+in_buf[600]*(0)+in_buf[601]*(2)+in_buf[602]*(4)+in_buf[603]*(11)+in_buf[604]*(1)+in_buf[605]*(-2)+in_buf[606]*(-7)+in_buf[607]*(11)+in_buf[608]*(0)+in_buf[609]*(8)+in_buf[610]*(1)+in_buf[611]*(3)+in_buf[612]*(9)+in_buf[613]*(32)+in_buf[614]*(23)+in_buf[615]*(-2)+in_buf[616]*(-21)+in_buf[617]*(-19)+in_buf[618]*(0)+in_buf[619]*(-33)+in_buf[620]*(-28)+in_buf[621]*(-21)+in_buf[622]*(-14)+in_buf[623]*(-2)+in_buf[624]*(10)+in_buf[625]*(19)+in_buf[626]*(11)+in_buf[627]*(4)+in_buf[628]*(-4)+in_buf[629]*(1)+in_buf[630]*(13)+in_buf[631]*(-2)+in_buf[632]*(-18)+in_buf[633]*(-14)+in_buf[634]*(-6)+in_buf[635]*(-3)+in_buf[636]*(-1)+in_buf[637]*(0)+in_buf[638]*(-7)+in_buf[639]*(12)+in_buf[640]*(19)+in_buf[641]*(23)+in_buf[642]*(-17)+in_buf[643]*(-3)+in_buf[644]*(4)+in_buf[645]*(4)+in_buf[646]*(-13)+in_buf[647]*(-42)+in_buf[648]*(-25)+in_buf[649]*(-14)+in_buf[650]*(5)+in_buf[651]*(18)+in_buf[652]*(15)+in_buf[653]*(21)+in_buf[654]*(5)+in_buf[655]*(9)+in_buf[656]*(19)+in_buf[657]*(17)+in_buf[658]*(10)+in_buf[659]*(3)+in_buf[660]*(0)+in_buf[661]*(-5)+in_buf[662]*(4)+in_buf[663]*(17)+in_buf[664]*(5)+in_buf[665]*(11)+in_buf[666]*(15)+in_buf[667]*(23)+in_buf[668]*(14)+in_buf[669]*(11)+in_buf[670]*(-22)+in_buf[671]*(-3)+in_buf[672]*(-3)+in_buf[673]*(-3)+in_buf[674]*(2)+in_buf[675]*(-27)+in_buf[676]*(-1)+in_buf[677]*(-7)+in_buf[678]*(0)+in_buf[679]*(-18)+in_buf[680]*(-10)+in_buf[681]*(-2)+in_buf[682]*(-13)+in_buf[683]*(-11)+in_buf[684]*(-8)+in_buf[685]*(0)+in_buf[686]*(7)+in_buf[687]*(17)+in_buf[688]*(-2)+in_buf[689]*(-8)+in_buf[690]*(18)+in_buf[691]*(44)+in_buf[692]*(24)+in_buf[693]*(13)+in_buf[694]*(16)+in_buf[695]*(24)+in_buf[696]*(53)+in_buf[697]*(4)+in_buf[698]*(7)+in_buf[699]*(-2)+in_buf[700]*(4)+in_buf[701]*(1)+in_buf[702]*(-13)+in_buf[703]*(14)+in_buf[704]*(15)+in_buf[705]*(-12)+in_buf[706]*(1)+in_buf[707]*(0)+in_buf[708]*(12)+in_buf[709]*(-4)+in_buf[710]*(-8)+in_buf[711]*(-18)+in_buf[712]*(-26)+in_buf[713]*(-23)+in_buf[714]*(7)+in_buf[715]*(4)+in_buf[716]*(-5)+in_buf[717]*(-2)+in_buf[718]*(12)+in_buf[719]*(-5)+in_buf[720]*(-9)+in_buf[721]*(-21)+in_buf[722]*(-28)+in_buf[723]*(-32)+in_buf[724]*(-18)+in_buf[725]*(-6)+in_buf[726]*(12)+in_buf[727]*(3)+in_buf[728]*(1)+in_buf[729]*(1)+in_buf[730]*(-1)+in_buf[731]*(1)+in_buf[732]*(-33)+in_buf[733]*(-35)+in_buf[734]*(-28)+in_buf[735]*(10)+in_buf[736]*(30)+in_buf[737]*(0)+in_buf[738]*(-11)+in_buf[739]*(-15)+in_buf[740]*(-8)+in_buf[741]*(4)+in_buf[742]*(10)+in_buf[743]*(2)+in_buf[744]*(-13)+in_buf[745]*(-17)+in_buf[746]*(7)+in_buf[747]*(30)+in_buf[748]*(17)+in_buf[749]*(-12)+in_buf[750]*(-11)+in_buf[751]*(-6)+in_buf[752]*(-29)+in_buf[753]*(11)+in_buf[754]*(1)+in_buf[755]*(-2)+in_buf[756]*(3)+in_buf[757]*(4)+in_buf[758]*(-3)+in_buf[759]*(-3)+in_buf[760]*(32)+in_buf[761]*(31)+in_buf[762]*(28)+in_buf[763]*(23)+in_buf[764]*(25)+in_buf[765]*(32)+in_buf[766]*(43)+in_buf[767]*(32)+in_buf[768]*(21)+in_buf[769]*(59)+in_buf[770]*(13)+in_buf[771]*(-4)+in_buf[772]*(8)+in_buf[773]*(40)+in_buf[774]*(21)+in_buf[775]*(12)+in_buf[776]*(1)+in_buf[777]*(-11)+in_buf[778]*(-2)+in_buf[779]*(7)+in_buf[780]*(3)+in_buf[781]*(3)+in_buf[782]*(3)+in_buf[783]*(-3);
assign in_buf_weight047=in_buf[0]*(0)+in_buf[1]*(-2)+in_buf[2]*(0)+in_buf[3]*(0)+in_buf[4]*(3)+in_buf[5]*(2)+in_buf[6]*(5)+in_buf[7]*(-4)+in_buf[8]*(2)+in_buf[9]*(-3)+in_buf[10]*(1)+in_buf[11]*(-2)+in_buf[12]*(3)+in_buf[13]*(-1)+in_buf[14]*(3)+in_buf[15]*(4)+in_buf[16]*(-3)+in_buf[17]*(4)+in_buf[18]*(-2)+in_buf[19]*(1)+in_buf[20]*(0)+in_buf[21]*(0)+in_buf[22]*(-3)+in_buf[23]*(1)+in_buf[24]*(2)+in_buf[25]*(3)+in_buf[26]*(2)+in_buf[27]*(2)+in_buf[28]*(1)+in_buf[29]*(-3)+in_buf[30]*(0)+in_buf[31]*(0)+in_buf[32]*(4)+in_buf[33]*(2)+in_buf[34]*(-2)+in_buf[35]*(0)+in_buf[36]*(-7)+in_buf[37]*(-2)+in_buf[38]*(0)+in_buf[39]*(3)+in_buf[40]*(-9)+in_buf[41]*(-7)+in_buf[42]*(-17)+in_buf[43]*(-15)+in_buf[44]*(-12)+in_buf[45]*(-1)+in_buf[46]*(0)+in_buf[47]*(-6)+in_buf[48]*(-9)+in_buf[49]*(-17)+in_buf[50]*(4)+in_buf[51]*(4)+in_buf[52]*(-3)+in_buf[53]*(2)+in_buf[54]*(0)+in_buf[55]*(-4)+in_buf[56]*(1)+in_buf[57]*(0)+in_buf[58]*(-3)+in_buf[59]*(0)+in_buf[60]*(0)+in_buf[61]*(-5)+in_buf[62]*(-2)+in_buf[63]*(-4)+in_buf[64]*(-13)+in_buf[65]*(4)+in_buf[66]*(19)+in_buf[67]*(7)+in_buf[68]*(-33)+in_buf[69]*(-23)+in_buf[70]*(22)+in_buf[71]*(48)+in_buf[72]*(34)+in_buf[73]*(21)+in_buf[74]*(24)+in_buf[75]*(11)+in_buf[76]*(17)+in_buf[77]*(2)+in_buf[78]*(15)+in_buf[79]*(22)+in_buf[80]*(3)+in_buf[81]*(-1)+in_buf[82]*(-3)+in_buf[83]*(1)+in_buf[84]*(-2)+in_buf[85]*(0)+in_buf[86]*(6)+in_buf[87]*(1)+in_buf[88]*(25)+in_buf[89]*(22)+in_buf[90]*(22)+in_buf[91]*(27)+in_buf[92]*(60)+in_buf[93]*(25)+in_buf[94]*(25)+in_buf[95]*(13)+in_buf[96]*(5)+in_buf[97]*(-9)+in_buf[98]*(-15)+in_buf[99]*(13)+in_buf[100]*(-10)+in_buf[101]*(-17)+in_buf[102]*(-7)+in_buf[103]*(-18)+in_buf[104]*(3)+in_buf[105]*(-12)+in_buf[106]*(-22)+in_buf[107]*(-13)+in_buf[108]*(28)+in_buf[109]*(-11)+in_buf[110]*(-3)+in_buf[111]*(2)+in_buf[112]*(1)+in_buf[113]*(6)+in_buf[114]*(6)+in_buf[115]*(25)+in_buf[116]*(22)+in_buf[117]*(18)+in_buf[118]*(25)+in_buf[119]*(49)+in_buf[120]*(43)+in_buf[121]*(26)+in_buf[122]*(34)+in_buf[123]*(39)+in_buf[124]*(21)+in_buf[125]*(10)+in_buf[126]*(7)+in_buf[127]*(22)+in_buf[128]*(13)+in_buf[129]*(8)+in_buf[130]*(29)+in_buf[131]*(21)+in_buf[132]*(1)+in_buf[133]*(-4)+in_buf[134]*(-10)+in_buf[135]*(-38)+in_buf[136]*(0)+in_buf[137]*(11)+in_buf[138]*(33)+in_buf[139]*(-1)+in_buf[140]*(-2)+in_buf[141]*(0)+in_buf[142]*(8)+in_buf[143]*(9)+in_buf[144]*(25)+in_buf[145]*(19)+in_buf[146]*(18)+in_buf[147]*(33)+in_buf[148]*(19)+in_buf[149]*(16)+in_buf[150]*(16)+in_buf[151]*(27)+in_buf[152]*(17)+in_buf[153]*(15)+in_buf[154]*(-2)+in_buf[155]*(8)+in_buf[156]*(11)+in_buf[157]*(15)+in_buf[158]*(16)+in_buf[159]*(8)+in_buf[160]*(7)+in_buf[161]*(-12)+in_buf[162]*(-20)+in_buf[163]*(-13)+in_buf[164]*(-12)+in_buf[165]*(-6)+in_buf[166]*(7)+in_buf[167]*(-1)+in_buf[168]*(-3)+in_buf[169]*(15)+in_buf[170]*(-17)+in_buf[171]*(-19)+in_buf[172]*(-5)+in_buf[173]*(5)+in_buf[174]*(3)+in_buf[175]*(2)+in_buf[176]*(13)+in_buf[177]*(10)+in_buf[178]*(9)+in_buf[179]*(9)+in_buf[180]*(0)+in_buf[181]*(10)+in_buf[182]*(8)+in_buf[183]*(6)+in_buf[184]*(23)+in_buf[185]*(10)+in_buf[186]*(4)+in_buf[187]*(4)+in_buf[188]*(-2)+in_buf[189]*(-13)+in_buf[190]*(-21)+in_buf[191]*(2)+in_buf[192]*(6)+in_buf[193]*(20)+in_buf[194]*(28)+in_buf[195]*(3)+in_buf[196]*(-1)+in_buf[197]*(23)+in_buf[198]*(-26)+in_buf[199]*(-11)+in_buf[200]*(9)+in_buf[201]*(26)+in_buf[202]*(3)+in_buf[203]*(-8)+in_buf[204]*(1)+in_buf[205]*(1)+in_buf[206]*(8)+in_buf[207]*(5)+in_buf[208]*(9)+in_buf[209]*(1)+in_buf[210]*(5)+in_buf[211]*(1)+in_buf[212]*(15)+in_buf[213]*(7)+in_buf[214]*(-9)+in_buf[215]*(8)+in_buf[216]*(18)+in_buf[217]*(8)+in_buf[218]*(-4)+in_buf[219]*(-8)+in_buf[220]*(1)+in_buf[221]*(33)+in_buf[222]*(-12)+in_buf[223]*(0)+in_buf[224]*(-2)+in_buf[225]*(-26)+in_buf[226]*(-17)+in_buf[227]*(14)+in_buf[228]*(13)+in_buf[229]*(22)+in_buf[230]*(-5)+in_buf[231]*(-9)+in_buf[232]*(7)+in_buf[233]*(10)+in_buf[234]*(18)+in_buf[235]*(10)+in_buf[236]*(-4)+in_buf[237]*(-6)+in_buf[238]*(-6)+in_buf[239]*(-6)+in_buf[240]*(6)+in_buf[241]*(-13)+in_buf[242]*(-6)+in_buf[243]*(-4)+in_buf[244]*(-1)+in_buf[245]*(14)+in_buf[246]*(14)+in_buf[247]*(-4)+in_buf[248]*(-8)+in_buf[249]*(13)+in_buf[250]*(-20)+in_buf[251]*(-7)+in_buf[252]*(-13)+in_buf[253]*(-23)+in_buf[254]*(11)+in_buf[255]*(6)+in_buf[256]*(0)+in_buf[257]*(10)+in_buf[258]*(9)+in_buf[259]*(3)+in_buf[260]*(19)+in_buf[261]*(12)+in_buf[262]*(13)+in_buf[263]*(3)+in_buf[264]*(-7)+in_buf[265]*(-12)+in_buf[266]*(-18)+in_buf[267]*(-12)+in_buf[268]*(-8)+in_buf[269]*(-17)+in_buf[270]*(-13)+in_buf[271]*(-19)+in_buf[272]*(-15)+in_buf[273]*(11)+in_buf[274]*(22)+in_buf[275]*(0)+in_buf[276]*(-36)+in_buf[277]*(0)+in_buf[278]*(-20)+in_buf[279]*(-3)+in_buf[280]*(-13)+in_buf[281]*(-15)+in_buf[282]*(-5)+in_buf[283]*(21)+in_buf[284]*(-3)+in_buf[285]*(-7)+in_buf[286]*(3)+in_buf[287]*(19)+in_buf[288]*(25)+in_buf[289]*(3)+in_buf[290]*(5)+in_buf[291]*(2)+in_buf[292]*(-2)+in_buf[293]*(-6)+in_buf[294]*(-7)+in_buf[295]*(-15)+in_buf[296]*(-13)+in_buf[297]*(-4)+in_buf[298]*(-4)+in_buf[299]*(-3)+in_buf[300]*(-1)+in_buf[301]*(1)+in_buf[302]*(2)+in_buf[303]*(-33)+in_buf[304]*(-59)+in_buf[305]*(6)+in_buf[306]*(15)+in_buf[307]*(9)+in_buf[308]*(-3)+in_buf[309]*(-31)+in_buf[310]*(-19)+in_buf[311]*(-2)+in_buf[312]*(-4)+in_buf[313]*(-23)+in_buf[314]*(-16)+in_buf[315]*(-6)+in_buf[316]*(8)+in_buf[317]*(-7)+in_buf[318]*(8)+in_buf[319]*(17)+in_buf[320]*(30)+in_buf[321]*(24)+in_buf[322]*(22)+in_buf[323]*(15)+in_buf[324]*(12)+in_buf[325]*(21)+in_buf[326]*(21)+in_buf[327]*(8)+in_buf[328]*(18)+in_buf[329]*(-4)+in_buf[330]*(-29)+in_buf[331]*(-62)+in_buf[332]*(-56)+in_buf[333]*(-4)+in_buf[334]*(-10)+in_buf[335]*(-5)+in_buf[336]*(0)+in_buf[337]*(-25)+in_buf[338]*(-5)+in_buf[339]*(-37)+in_buf[340]*(-38)+in_buf[341]*(-27)+in_buf[342]*(-25)+in_buf[343]*(-10)+in_buf[344]*(4)+in_buf[345]*(7)+in_buf[346]*(23)+in_buf[347]*(29)+in_buf[348]*(29)+in_buf[349]*(34)+in_buf[350]*(27)+in_buf[351]*(21)+in_buf[352]*(14)+in_buf[353]*(11)+in_buf[354]*(19)+in_buf[355]*(19)+in_buf[356]*(11)+in_buf[357]*(0)+in_buf[358]*(-12)+in_buf[359]*(-31)+in_buf[360]*(-73)+in_buf[361]*(-30)+in_buf[362]*(20)+in_buf[363]*(-6)+in_buf[364]*(20)+in_buf[365]*(-11)+in_buf[366]*(-26)+in_buf[367]*(-52)+in_buf[368]*(-41)+in_buf[369]*(-34)+in_buf[370]*(-29)+in_buf[371]*(-7)+in_buf[372]*(-3)+in_buf[373]*(0)+in_buf[374]*(7)+in_buf[375]*(18)+in_buf[376]*(33)+in_buf[377]*(34)+in_buf[378]*(33)+in_buf[379]*(15)+in_buf[380]*(20)+in_buf[381]*(2)+in_buf[382]*(5)+in_buf[383]*(0)+in_buf[384]*(-3)+in_buf[385]*(0)+in_buf[386]*(-1)+in_buf[387]*(-11)+in_buf[388]*(-1)+in_buf[389]*(-34)+in_buf[390]*(-3)+in_buf[391]*(-14)+in_buf[392]*(-12)+in_buf[393]*(0)+in_buf[394]*(-24)+in_buf[395]*(-38)+in_buf[396]*(-55)+in_buf[397]*(-76)+in_buf[398]*(-47)+in_buf[399]*(-13)+in_buf[400]*(-23)+in_buf[401]*(-19)+in_buf[402]*(0)+in_buf[403]*(10)+in_buf[404]*(33)+in_buf[405]*(40)+in_buf[406]*(33)+in_buf[407]*(14)+in_buf[408]*(4)+in_buf[409]*(8)+in_buf[410]*(-1)+in_buf[411]*(-17)+in_buf[412]*(-2)+in_buf[413]*(2)+in_buf[414]*(1)+in_buf[415]*(9)+in_buf[416]*(37)+in_buf[417]*(-17)+in_buf[418]*(-3)+in_buf[419]*(-18)+in_buf[420]*(-15)+in_buf[421]*(11)+in_buf[422]*(20)+in_buf[423]*(-19)+in_buf[424]*(-37)+in_buf[425]*(-86)+in_buf[426]*(-66)+in_buf[427]*(-68)+in_buf[428]*(-57)+in_buf[429]*(-49)+in_buf[430]*(-20)+in_buf[431]*(-4)+in_buf[432]*(16)+in_buf[433]*(22)+in_buf[434]*(10)+in_buf[435]*(-7)+in_buf[436]*(-8)+in_buf[437]*(0)+in_buf[438]*(0)+in_buf[439]*(-4)+in_buf[440]*(3)+in_buf[441]*(20)+in_buf[442]*(29)+in_buf[443]*(41)+in_buf[444]*(44)+in_buf[445]*(11)+in_buf[446]*(22)+in_buf[447]*(-19)+in_buf[448]*(-3)+in_buf[449]*(18)+in_buf[450]*(31)+in_buf[451]*(4)+in_buf[452]*(-10)+in_buf[453]*(-53)+in_buf[454]*(-58)+in_buf[455]*(-73)+in_buf[456]*(-79)+in_buf[457]*(-79)+in_buf[458]*(-74)+in_buf[459]*(-71)+in_buf[460]*(-50)+in_buf[461]*(-24)+in_buf[462]*(-24)+in_buf[463]*(-18)+in_buf[464]*(-2)+in_buf[465]*(4)+in_buf[466]*(29)+in_buf[467]*(8)+in_buf[468]*(0)+in_buf[469]*(7)+in_buf[470]*(33)+in_buf[471]*(39)+in_buf[472]*(40)+in_buf[473]*(22)+in_buf[474]*(-3)+in_buf[475]*(-17)+in_buf[476]*(-4)+in_buf[477]*(14)+in_buf[478]*(20)+in_buf[479]*(11)+in_buf[480]*(-10)+in_buf[481]*(-11)+in_buf[482]*(-20)+in_buf[483]*(-48)+in_buf[484]*(-54)+in_buf[485]*(-78)+in_buf[486]*(-90)+in_buf[487]*(-115)+in_buf[488]*(-114)+in_buf[489]*(-72)+in_buf[490]*(-46)+in_buf[491]*(-13)+in_buf[492]*(-5)+in_buf[493]*(13)+in_buf[494]*(14)+in_buf[495]*(15)+in_buf[496]*(8)+in_buf[497]*(10)+in_buf[498]*(8)+in_buf[499]*(28)+in_buf[500]*(7)+in_buf[501]*(-36)+in_buf[502]*(-5)+in_buf[503]*(-7)+in_buf[504]*(-16)+in_buf[505]*(8)+in_buf[506]*(3)+in_buf[507]*(41)+in_buf[508]*(16)+in_buf[509]*(25)+in_buf[510]*(21)+in_buf[511]*(-25)+in_buf[512]*(-31)+in_buf[513]*(-29)+in_buf[514]*(-41)+in_buf[515]*(-49)+in_buf[516]*(-79)+in_buf[517]*(-44)+in_buf[518]*(-22)+in_buf[519]*(-13)+in_buf[520]*(7)+in_buf[521]*(8)+in_buf[522]*(7)+in_buf[523]*(22)+in_buf[524]*(10)+in_buf[525]*(7)+in_buf[526]*(9)+in_buf[527]*(23)+in_buf[528]*(33)+in_buf[529]*(7)+in_buf[530]*(-35)+in_buf[531]*(-17)+in_buf[532]*(7)+in_buf[533]*(-36)+in_buf[534]*(-23)+in_buf[535]*(33)+in_buf[536]*(24)+in_buf[537]*(35)+in_buf[538]*(40)+in_buf[539]*(13)+in_buf[540]*(-8)+in_buf[541]*(0)+in_buf[542]*(7)+in_buf[543]*(16)+in_buf[544]*(-6)+in_buf[545]*(-6)+in_buf[546]*(-7)+in_buf[547]*(-8)+in_buf[548]*(5)+in_buf[549]*(-5)+in_buf[550]*(9)+in_buf[551]*(10)+in_buf[552]*(5)+in_buf[553]*(11)+in_buf[554]*(0)+in_buf[555]*(32)+in_buf[556]*(38)+in_buf[557]*(23)+in_buf[558]*(-45)+in_buf[559]*(-21)+in_buf[560]*(0)+in_buf[561]*(13)+in_buf[562]*(-27)+in_buf[563]*(20)+in_buf[564]*(31)+in_buf[565]*(31)+in_buf[566]*(33)+in_buf[567]*(15)+in_buf[568]*(12)+in_buf[569]*(18)+in_buf[570]*(15)+in_buf[571]*(23)+in_buf[572]*(4)+in_buf[573]*(6)+in_buf[574]*(4)+in_buf[575]*(-9)+in_buf[576]*(-5)+in_buf[577]*(-2)+in_buf[578]*(8)+in_buf[579]*(4)+in_buf[580]*(11)+in_buf[581]*(11)+in_buf[582]*(17)+in_buf[583]*(17)+in_buf[584]*(13)+in_buf[585]*(-36)+in_buf[586]*(-31)+in_buf[587]*(2)+in_buf[588]*(0)+in_buf[589]*(15)+in_buf[590]*(-13)+in_buf[591]*(-6)+in_buf[592]*(24)+in_buf[593]*(22)+in_buf[594]*(22)+in_buf[595]*(23)+in_buf[596]*(35)+in_buf[597]*(26)+in_buf[598]*(25)+in_buf[599]*(22)+in_buf[600]*(17)+in_buf[601]*(8)+in_buf[602]*(-1)+in_buf[603]*(-4)+in_buf[604]*(-4)+in_buf[605]*(-6)+in_buf[606]*(-2)+in_buf[607]*(3)+in_buf[608]*(15)+in_buf[609]*(-4)+in_buf[610]*(-17)+in_buf[611]*(14)+in_buf[612]*(-38)+in_buf[613]*(-44)+in_buf[614]*(-21)+in_buf[615]*(-1)+in_buf[616]*(-1)+in_buf[617]*(27)+in_buf[618]*(-9)+in_buf[619]*(11)+in_buf[620]*(14)+in_buf[621]*(6)+in_buf[622]*(-7)+in_buf[623]*(3)+in_buf[624]*(18)+in_buf[625]*(13)+in_buf[626]*(21)+in_buf[627]*(7)+in_buf[628]*(2)+in_buf[629]*(0)+in_buf[630]*(2)+in_buf[631]*(-1)+in_buf[632]*(8)+in_buf[633]*(6)+in_buf[634]*(0)+in_buf[635]*(-2)+in_buf[636]*(2)+in_buf[637]*(-15)+in_buf[638]*(18)+in_buf[639]*(10)+in_buf[640]*(-52)+in_buf[641]*(-29)+in_buf[642]*(11)+in_buf[643]*(-2)+in_buf[644]*(-1)+in_buf[645]*(5)+in_buf[646]*(27)+in_buf[647]*(50)+in_buf[648]*(40)+in_buf[649]*(23)+in_buf[650]*(-3)+in_buf[651]*(-7)+in_buf[652]*(2)+in_buf[653]*(0)+in_buf[654]*(7)+in_buf[655]*(17)+in_buf[656]*(8)+in_buf[657]*(18)+in_buf[658]*(8)+in_buf[659]*(8)+in_buf[660]*(8)+in_buf[661]*(2)+in_buf[662]*(2)+in_buf[663]*(-10)+in_buf[664]*(-4)+in_buf[665]*(-12)+in_buf[666]*(-14)+in_buf[667]*(-15)+in_buf[668]*(-34)+in_buf[669]*(-19)+in_buf[670]*(22)+in_buf[671]*(1)+in_buf[672]*(-1)+in_buf[673]*(-1)+in_buf[674]*(0)+in_buf[675]*(32)+in_buf[676]*(48)+in_buf[677]*(27)+in_buf[678]*(6)+in_buf[679]*(27)+in_buf[680]*(9)+in_buf[681]*(-14)+in_buf[682]*(-1)+in_buf[683]*(-4)+in_buf[684]*(-5)+in_buf[685]*(-5)+in_buf[686]*(-11)+in_buf[687]*(-1)+in_buf[688]*(6)+in_buf[689]*(-9)+in_buf[690]*(-22)+in_buf[691]*(-46)+in_buf[692]*(-33)+in_buf[693]*(-32)+in_buf[694]*(-25)+in_buf[695]*(10)+in_buf[696]*(-21)+in_buf[697]*(1)+in_buf[698]*(0)+in_buf[699]*(1)+in_buf[700]*(-3)+in_buf[701]*(4)+in_buf[702]*(7)+in_buf[703]*(-9)+in_buf[704]*(24)+in_buf[705]*(23)+in_buf[706]*(7)+in_buf[707]*(24)+in_buf[708]*(14)+in_buf[709]*(11)+in_buf[710]*(33)+in_buf[711]*(0)+in_buf[712]*(21)+in_buf[713]*(24)+in_buf[714]*(4)+in_buf[715]*(-4)+in_buf[716]*(-12)+in_buf[717]*(-17)+in_buf[718]*(-24)+in_buf[719]*(-36)+in_buf[720]*(-15)+in_buf[721]*(-24)+in_buf[722]*(-13)+in_buf[723]*(2)+in_buf[724]*(7)+in_buf[725]*(7)+in_buf[726]*(-1)+in_buf[727]*(-3)+in_buf[728]*(-1)+in_buf[729]*(0)+in_buf[730]*(4)+in_buf[731]*(11)+in_buf[732]*(26)+in_buf[733]*(28)+in_buf[734]*(8)+in_buf[735]*(-3)+in_buf[736]*(-17)+in_buf[737]*(15)+in_buf[738]*(26)+in_buf[739]*(10)+in_buf[740]*(-5)+in_buf[741]*(0)+in_buf[742]*(19)+in_buf[743]*(12)+in_buf[744]*(4)+in_buf[745]*(11)+in_buf[746]*(21)+in_buf[747]*(-5)+in_buf[748]*(-1)+in_buf[749]*(5)+in_buf[750]*(-9)+in_buf[751]*(-8)+in_buf[752]*(0)+in_buf[753]*(1)+in_buf[754]*(-3)+in_buf[755]*(0)+in_buf[756]*(-2)+in_buf[757]*(4)+in_buf[758]*(-1)+in_buf[759]*(0)+in_buf[760]*(-4)+in_buf[761]*(-5)+in_buf[762]*(-26)+in_buf[763]*(-26)+in_buf[764]*(-27)+in_buf[765]*(-26)+in_buf[766]*(-33)+in_buf[767]*(-32)+in_buf[768]*(-43)+in_buf[769]*(-10)+in_buf[770]*(-2)+in_buf[771]*(15)+in_buf[772]*(-3)+in_buf[773]*(-35)+in_buf[774]*(-32)+in_buf[775]*(-38)+in_buf[776]*(-24)+in_buf[777]*(3)+in_buf[778]*(-2)+in_buf[779]*(-3)+in_buf[780]*(-2)+in_buf[781]*(1)+in_buf[782]*(1)+in_buf[783]*(-3);
assign in_buf_weight048=in_buf[0]*(0)+in_buf[1]*(3)+in_buf[2]*(2)+in_buf[3]*(-1)+in_buf[4]*(-3)+in_buf[5]*(0)+in_buf[6]*(-2)+in_buf[7]*(4)+in_buf[8]*(-2)+in_buf[9]*(0)+in_buf[10]*(0)+in_buf[11]*(3)+in_buf[12]*(15)+in_buf[13]*(13)+in_buf[14]*(-4)+in_buf[15]*(-5)+in_buf[16]*(3)+in_buf[17]*(3)+in_buf[18]*(5)+in_buf[19]*(2)+in_buf[20]*(0)+in_buf[21]*(-2)+in_buf[22]*(-1)+in_buf[23]*(4)+in_buf[24]*(-2)+in_buf[25]*(-3)+in_buf[26]*(1)+in_buf[27]*(0)+in_buf[28]*(0)+in_buf[29]*(1)+in_buf[30]*(1)+in_buf[31]*(2)+in_buf[32]*(7)+in_buf[33]*(5)+in_buf[34]*(8)+in_buf[35]*(9)+in_buf[36]*(17)+in_buf[37]*(12)+in_buf[38]*(18)+in_buf[39]*(5)+in_buf[40]*(10)+in_buf[41]*(0)+in_buf[42]*(-10)+in_buf[43]*(38)+in_buf[44]*(14)+in_buf[45]*(27)+in_buf[46]*(34)+in_buf[47]*(32)+in_buf[48]*(24)+in_buf[49]*(22)+in_buf[50]*(15)+in_buf[51]*(14)+in_buf[52]*(4)+in_buf[53]*(1)+in_buf[54]*(4)+in_buf[55]*(-2)+in_buf[56]*(-1)+in_buf[57]*(3)+in_buf[58]*(16)+in_buf[59]*(21)+in_buf[60]*(34)+in_buf[61]*(4)+in_buf[62]*(18)+in_buf[63]*(17)+in_buf[64]*(4)+in_buf[65]*(4)+in_buf[66]*(16)+in_buf[67]*(29)+in_buf[68]*(40)+in_buf[69]*(42)+in_buf[70]*(17)+in_buf[71]*(4)+in_buf[72]*(-3)+in_buf[73]*(12)+in_buf[74]*(45)+in_buf[75]*(41)+in_buf[76]*(34)+in_buf[77]*(32)+in_buf[78]*(40)+in_buf[79]*(5)+in_buf[80]*(-2)+in_buf[81]*(-2)+in_buf[82]*(2)+in_buf[83]*(-1)+in_buf[84]*(0)+in_buf[85]*(-3)+in_buf[86]*(19)+in_buf[87]*(24)+in_buf[88]*(15)+in_buf[89]*(-14)+in_buf[90]*(25)+in_buf[91]*(-12)+in_buf[92]*(-37)+in_buf[93]*(-22)+in_buf[94]*(-7)+in_buf[95]*(-6)+in_buf[96]*(-7)+in_buf[97]*(0)+in_buf[98]*(-9)+in_buf[99]*(-1)+in_buf[100]*(7)+in_buf[101]*(0)+in_buf[102]*(5)+in_buf[103]*(10)+in_buf[104]*(9)+in_buf[105]*(37)+in_buf[106]*(31)+in_buf[107]*(21)+in_buf[108]*(-3)+in_buf[109]*(-14)+in_buf[110]*(-22)+in_buf[111]*(-1)+in_buf[112]*(4)+in_buf[113]*(-1)+in_buf[114]*(0)+in_buf[115]*(-22)+in_buf[116]*(-8)+in_buf[117]*(-2)+in_buf[118]*(-26)+in_buf[119]*(-19)+in_buf[120]*(-3)+in_buf[121]*(-4)+in_buf[122]*(3)+in_buf[123]*(0)+in_buf[124]*(13)+in_buf[125]*(12)+in_buf[126]*(19)+in_buf[127]*(17)+in_buf[128]*(15)+in_buf[129]*(-3)+in_buf[130]*(-23)+in_buf[131]*(-8)+in_buf[132]*(-14)+in_buf[133]*(2)+in_buf[134]*(2)+in_buf[135]*(0)+in_buf[136]*(3)+in_buf[137]*(-20)+in_buf[138]*(31)+in_buf[139]*(17)+in_buf[140]*(-1)+in_buf[141]*(1)+in_buf[142]*(13)+in_buf[143]*(-23)+in_buf[144]*(2)+in_buf[145]*(5)+in_buf[146]*(1)+in_buf[147]*(1)+in_buf[148]*(-10)+in_buf[149]*(-1)+in_buf[150]*(-9)+in_buf[151]*(16)+in_buf[152]*(24)+in_buf[153]*(21)+in_buf[154]*(16)+in_buf[155]*(10)+in_buf[156]*(0)+in_buf[157]*(-1)+in_buf[158]*(-6)+in_buf[159]*(0)+in_buf[160]*(-2)+in_buf[161]*(0)+in_buf[162]*(-12)+in_buf[163]*(-27)+in_buf[164]*(6)+in_buf[165]*(21)+in_buf[166]*(21)+in_buf[167]*(5)+in_buf[168]*(1)+in_buf[169]*(-15)+in_buf[170]*(-25)+in_buf[171]*(-10)+in_buf[172]*(-25)+in_buf[173]*(-32)+in_buf[174]*(-13)+in_buf[175]*(-8)+in_buf[176]*(-7)+in_buf[177]*(6)+in_buf[178]*(8)+in_buf[179]*(21)+in_buf[180]*(16)+in_buf[181]*(11)+in_buf[182]*(18)+in_buf[183]*(5)+in_buf[184]*(8)+in_buf[185]*(16)+in_buf[186]*(1)+in_buf[187]*(-10)+in_buf[188]*(-6)+in_buf[189]*(-4)+in_buf[190]*(-13)+in_buf[191]*(-16)+in_buf[192]*(-18)+in_buf[193]*(40)+in_buf[194]*(10)+in_buf[195]*(-10)+in_buf[196]*(2)+in_buf[197]*(-22)+in_buf[198]*(-12)+in_buf[199]*(-9)+in_buf[200]*(-40)+in_buf[201]*(-54)+in_buf[202]*(-5)+in_buf[203]*(-4)+in_buf[204]*(-1)+in_buf[205]*(10)+in_buf[206]*(15)+in_buf[207]*(1)+in_buf[208]*(1)+in_buf[209]*(-1)+in_buf[210]*(-13)+in_buf[211]*(3)+in_buf[212]*(3)+in_buf[213]*(-6)+in_buf[214]*(0)+in_buf[215]*(-4)+in_buf[216]*(-3)+in_buf[217]*(0)+in_buf[218]*(2)+in_buf[219]*(-1)+in_buf[220]*(0)+in_buf[221]*(18)+in_buf[222]*(-13)+in_buf[223]*(-26)+in_buf[224]*(-14)+in_buf[225]*(15)+in_buf[226]*(-14)+in_buf[227]*(13)+in_buf[228]*(-12)+in_buf[229]*(-4)+in_buf[230]*(18)+in_buf[231]*(11)+in_buf[232]*(23)+in_buf[233]*(4)+in_buf[234]*(8)+in_buf[235]*(-8)+in_buf[236]*(-15)+in_buf[237]*(-15)+in_buf[238]*(-6)+in_buf[239]*(-3)+in_buf[240]*(-4)+in_buf[241]*(-4)+in_buf[242]*(-4)+in_buf[243]*(10)+in_buf[244]*(-4)+in_buf[245]*(0)+in_buf[246]*(-6)+in_buf[247]*(-2)+in_buf[248]*(-9)+in_buf[249]*(7)+in_buf[250]*(18)+in_buf[251]*(14)+in_buf[252]*(9)+in_buf[253]*(17)+in_buf[254]*(-10)+in_buf[255]*(18)+in_buf[256]*(-14)+in_buf[257]*(-1)+in_buf[258]*(15)+in_buf[259]*(6)+in_buf[260]*(8)+in_buf[261]*(7)+in_buf[262]*(4)+in_buf[263]*(-4)+in_buf[264]*(-13)+in_buf[265]*(2)+in_buf[266]*(5)+in_buf[267]*(3)+in_buf[268]*(-6)+in_buf[269]*(-4)+in_buf[270]*(-10)+in_buf[271]*(3)+in_buf[272]*(10)+in_buf[273]*(10)+in_buf[274]*(2)+in_buf[275]*(-1)+in_buf[276]*(-19)+in_buf[277]*(14)+in_buf[278]*(16)+in_buf[279]*(17)+in_buf[280]*(9)+in_buf[281]*(3)+in_buf[282]*(-19)+in_buf[283]*(-11)+in_buf[284]*(3)+in_buf[285]*(2)+in_buf[286]*(21)+in_buf[287]*(12)+in_buf[288]*(0)+in_buf[289]*(8)+in_buf[290]*(7)+in_buf[291]*(-4)+in_buf[292]*(3)+in_buf[293]*(11)+in_buf[294]*(33)+in_buf[295]*(14)+in_buf[296]*(-3)+in_buf[297]*(-18)+in_buf[298]*(-12)+in_buf[299]*(-1)+in_buf[300]*(13)+in_buf[301]*(11)+in_buf[302]*(4)+in_buf[303]*(23)+in_buf[304]*(-7)+in_buf[305]*(-7)+in_buf[306]*(-11)+in_buf[307]*(31)+in_buf[308]*(12)+in_buf[309]*(-12)+in_buf[310]*(30)+in_buf[311]*(26)+in_buf[312]*(21)+in_buf[313]*(25)+in_buf[314]*(15)+in_buf[315]*(20)+in_buf[316]*(14)+in_buf[317]*(14)+in_buf[318]*(-2)+in_buf[319]*(9)+in_buf[320]*(21)+in_buf[321]*(34)+in_buf[322]*(44)+in_buf[323]*(11)+in_buf[324]*(-1)+in_buf[325]*(-7)+in_buf[326]*(-1)+in_buf[327]*(5)+in_buf[328]*(25)+in_buf[329]*(19)+in_buf[330]*(14)+in_buf[331]*(13)+in_buf[332]*(17)+in_buf[333]*(5)+in_buf[334]*(12)+in_buf[335]*(19)+in_buf[336]*(14)+in_buf[337]*(4)+in_buf[338]*(31)+in_buf[339]*(59)+in_buf[340]*(34)+in_buf[341]*(17)+in_buf[342]*(18)+in_buf[343]*(17)+in_buf[344]*(13)+in_buf[345]*(9)+in_buf[346]*(-14)+in_buf[347]*(2)+in_buf[348]*(2)+in_buf[349]*(18)+in_buf[350]*(23)+in_buf[351]*(18)+in_buf[352]*(15)+in_buf[353]*(19)+in_buf[354]*(3)+in_buf[355]*(26)+in_buf[356]*(28)+in_buf[357]*(21)+in_buf[358]*(10)+in_buf[359]*(15)+in_buf[360]*(19)+in_buf[361]*(-1)+in_buf[362]*(13)+in_buf[363]*(35)+in_buf[364]*(8)+in_buf[365]*(-5)+in_buf[366]*(20)+in_buf[367]*(61)+in_buf[368]*(18)+in_buf[369]*(16)+in_buf[370]*(5)+in_buf[371]*(11)+in_buf[372]*(14)+in_buf[373]*(2)+in_buf[374]*(-12)+in_buf[375]*(4)+in_buf[376]*(2)+in_buf[377]*(11)+in_buf[378]*(20)+in_buf[379]*(27)+in_buf[380]*(21)+in_buf[381]*(10)+in_buf[382]*(14)+in_buf[383]*(20)+in_buf[384]*(33)+in_buf[385]*(13)+in_buf[386]*(25)+in_buf[387]*(14)+in_buf[388]*(-4)+in_buf[389]*(6)+in_buf[390]*(0)+in_buf[391]*(2)+in_buf[392]*(-17)+in_buf[393]*(-1)+in_buf[394]*(1)+in_buf[395]*(36)+in_buf[396]*(1)+in_buf[397]*(0)+in_buf[398]*(14)+in_buf[399]*(-4)+in_buf[400]*(0)+in_buf[401]*(-5)+in_buf[402]*(-4)+in_buf[403]*(8)+in_buf[404]*(6)+in_buf[405]*(14)+in_buf[406]*(19)+in_buf[407]*(13)+in_buf[408]*(19)+in_buf[409]*(9)+in_buf[410]*(16)+in_buf[411]*(19)+in_buf[412]*(10)+in_buf[413]*(1)+in_buf[414]*(2)+in_buf[415]*(10)+in_buf[416]*(-25)+in_buf[417]*(-5)+in_buf[418]*(-34)+in_buf[419]*(-3)+in_buf[420]*(-13)+in_buf[421]*(1)+in_buf[422]*(-22)+in_buf[423]*(7)+in_buf[424]*(-10)+in_buf[425]*(-6)+in_buf[426]*(-2)+in_buf[427]*(3)+in_buf[428]*(7)+in_buf[429]*(3)+in_buf[430]*(0)+in_buf[431]*(8)+in_buf[432]*(0)+in_buf[433]*(17)+in_buf[434]*(26)+in_buf[435]*(11)+in_buf[436]*(12)+in_buf[437]*(10)+in_buf[438]*(8)+in_buf[439]*(7)+in_buf[440]*(4)+in_buf[441]*(-8)+in_buf[442]*(-16)+in_buf[443]*(-28)+in_buf[444]*(-28)+in_buf[445]*(-10)+in_buf[446]*(-49)+in_buf[447]*(-16)+in_buf[448]*(5)+in_buf[449]*(1)+in_buf[450]*(-10)+in_buf[451]*(-22)+in_buf[452]*(-18)+in_buf[453]*(-3)+in_buf[454]*(8)+in_buf[455]*(-3)+in_buf[456]*(5)+in_buf[457]*(2)+in_buf[458]*(3)+in_buf[459]*(1)+in_buf[460]*(-3)+in_buf[461]*(-4)+in_buf[462]*(16)+in_buf[463]*(0)+in_buf[464]*(6)+in_buf[465]*(8)+in_buf[466]*(-11)+in_buf[467]*(-22)+in_buf[468]*(-10)+in_buf[469]*(-6)+in_buf[470]*(-17)+in_buf[471]*(-24)+in_buf[472]*(-22)+in_buf[473]*(-19)+in_buf[474]*(-51)+in_buf[475]*(-26)+in_buf[476]*(-1)+in_buf[477]*(0)+in_buf[478]*(-10)+in_buf[479]*(-43)+in_buf[480]*(-19)+in_buf[481]*(0)+in_buf[482]*(-8)+in_buf[483]*(-17)+in_buf[484]*(4)+in_buf[485]*(6)+in_buf[486]*(0)+in_buf[487]*(-1)+in_buf[488]*(-5)+in_buf[489]*(-7)+in_buf[490]*(6)+in_buf[491]*(-4)+in_buf[492]*(-5)+in_buf[493]*(-1)+in_buf[494]*(-13)+in_buf[495]*(-21)+in_buf[496]*(-6)+in_buf[497]*(-9)+in_buf[498]*(0)+in_buf[499]*(-10)+in_buf[500]*(5)+in_buf[501]*(-8)+in_buf[502]*(-25)+in_buf[503]*(-5)+in_buf[504]*(40)+in_buf[505]*(-4)+in_buf[506]*(8)+in_buf[507]*(-48)+in_buf[508]*(-21)+in_buf[509]*(-2)+in_buf[510]*(-9)+in_buf[511]*(-4)+in_buf[512]*(-2)+in_buf[513]*(0)+in_buf[514]*(0)+in_buf[515]*(-12)+in_buf[516]*(-20)+in_buf[517]*(-12)+in_buf[518]*(-10)+in_buf[519]*(-13)+in_buf[520]*(-18)+in_buf[521]*(-4)+in_buf[522]*(-10)+in_buf[523]*(-10)+in_buf[524]*(1)+in_buf[525]*(-10)+in_buf[526]*(1)+in_buf[527]*(4)+in_buf[528]*(0)+in_buf[529]*(10)+in_buf[530]*(-9)+in_buf[531]*(-17)+in_buf[532]*(8)+in_buf[533]*(33)+in_buf[534]*(2)+in_buf[535]*(-61)+in_buf[536]*(-15)+in_buf[537]*(-3)+in_buf[538]*(-5)+in_buf[539]*(-9)+in_buf[540]*(-1)+in_buf[541]*(0)+in_buf[542]*(0)+in_buf[543]*(-32)+in_buf[544]*(-26)+in_buf[545]*(-16)+in_buf[546]*(-19)+in_buf[547]*(-5)+in_buf[548]*(-5)+in_buf[549]*(-7)+in_buf[550]*(-12)+in_buf[551]*(-1)+in_buf[552]*(-4)+in_buf[553]*(-11)+in_buf[554]*(9)+in_buf[555]*(16)+in_buf[556]*(6)+in_buf[557]*(13)+in_buf[558]*(-45)+in_buf[559]*(-21)+in_buf[560]*(-3)+in_buf[561]*(8)+in_buf[562]*(0)+in_buf[563]*(-50)+in_buf[564]*(-8)+in_buf[565]*(0)+in_buf[566]*(-7)+in_buf[567]*(0)+in_buf[568]*(0)+in_buf[569]*(-9)+in_buf[570]*(-1)+in_buf[571]*(-11)+in_buf[572]*(-9)+in_buf[573]*(-9)+in_buf[574]*(-4)+in_buf[575]*(-1)+in_buf[576]*(-3)+in_buf[577]*(-15)+in_buf[578]*(-11)+in_buf[579]*(-4)+in_buf[580]*(1)+in_buf[581]*(1)+in_buf[582]*(9)+in_buf[583]*(2)+in_buf[584]*(19)+in_buf[585]*(5)+in_buf[586]*(-37)+in_buf[587]*(14)+in_buf[588]*(-9)+in_buf[589]*(-5)+in_buf[590]*(3)+in_buf[591]*(-13)+in_buf[592]*(2)+in_buf[593]*(0)+in_buf[594]*(17)+in_buf[595]*(9)+in_buf[596]*(2)+in_buf[597]*(4)+in_buf[598]*(5)+in_buf[599]*(5)+in_buf[600]*(8)+in_buf[601]*(4)+in_buf[602]*(-2)+in_buf[603]*(-3)+in_buf[604]*(0)+in_buf[605]*(-2)+in_buf[606]*(-6)+in_buf[607]*(0)+in_buf[608]*(2)+in_buf[609]*(-1)+in_buf[610]*(-5)+in_buf[611]*(-13)+in_buf[612]*(-26)+in_buf[613]*(-11)+in_buf[614]*(-34)+in_buf[615]*(1)+in_buf[616]*(-2)+in_buf[617]*(-9)+in_buf[618]*(-13)+in_buf[619]*(-6)+in_buf[620]*(18)+in_buf[621]*(9)+in_buf[622]*(17)+in_buf[623]*(19)+in_buf[624]*(10)+in_buf[625]*(12)+in_buf[626]*(9)+in_buf[627]*(3)+in_buf[628]*(5)+in_buf[629]*(3)+in_buf[630]*(-1)+in_buf[631]*(-4)+in_buf[632]*(-12)+in_buf[633]*(-11)+in_buf[634]*(-12)+in_buf[635]*(-23)+in_buf[636]*(-7)+in_buf[637]*(-14)+in_buf[638]*(-13)+in_buf[639]*(-19)+in_buf[640]*(-28)+in_buf[641]*(6)+in_buf[642]*(-19)+in_buf[643]*(0)+in_buf[644]*(-1)+in_buf[645]*(-3)+in_buf[646]*(-28)+in_buf[647]*(-32)+in_buf[648]*(-3)+in_buf[649]*(-2)+in_buf[650]*(-13)+in_buf[651]*(3)+in_buf[652]*(3)+in_buf[653]*(8)+in_buf[654]*(-9)+in_buf[655]*(-20)+in_buf[656]*(6)+in_buf[657]*(1)+in_buf[658]*(-9)+in_buf[659]*(-6)+in_buf[660]*(-7)+in_buf[661]*(-9)+in_buf[662]*(-9)+in_buf[663]*(-8)+in_buf[664]*(-9)+in_buf[665]*(-19)+in_buf[666]*(-4)+in_buf[667]*(0)+in_buf[668]*(-25)+in_buf[669]*(-14)+in_buf[670]*(-27)+in_buf[671]*(0)+in_buf[672]*(2)+in_buf[673]*(0)+in_buf[674]*(-8)+in_buf[675]*(-36)+in_buf[676]*(-28)+in_buf[677]*(6)+in_buf[678]*(0)+in_buf[679]*(6)+in_buf[680]*(0)+in_buf[681]*(-14)+in_buf[682]*(4)+in_buf[683]*(-8)+in_buf[684]*(-3)+in_buf[685]*(-8)+in_buf[686]*(-25)+in_buf[687]*(-11)+in_buf[688]*(-24)+in_buf[689]*(-40)+in_buf[690]*(-11)+in_buf[691]*(22)+in_buf[692]*(-7)+in_buf[693]*(-28)+in_buf[694]*(-25)+in_buf[695]*(-6)+in_buf[696]*(-21)+in_buf[697]*(-5)+in_buf[698]*(-11)+in_buf[699]*(0)+in_buf[700]*(-1)+in_buf[701]*(0)+in_buf[702]*(-6)+in_buf[703]*(-1)+in_buf[704]*(-30)+in_buf[705]*(-14)+in_buf[706]*(0)+in_buf[707]*(1)+in_buf[708]*(14)+in_buf[709]*(17)+in_buf[710]*(8)+in_buf[711]*(-2)+in_buf[712]*(0)+in_buf[713]*(-3)+in_buf[714]*(7)+in_buf[715]*(-12)+in_buf[716]*(-25)+in_buf[717]*(5)+in_buf[718]*(23)+in_buf[719]*(32)+in_buf[720]*(14)+in_buf[721]*(0)+in_buf[722]*(-21)+in_buf[723]*(-20)+in_buf[724]*(-8)+in_buf[725]*(0)+in_buf[726]*(-4)+in_buf[727]*(3)+in_buf[728]*(-1)+in_buf[729]*(-2)+in_buf[730]*(1)+in_buf[731]*(27)+in_buf[732]*(-3)+in_buf[733]*(0)+in_buf[734]*(17)+in_buf[735]*(28)+in_buf[736]*(35)+in_buf[737]*(48)+in_buf[738]*(32)+in_buf[739]*(16)+in_buf[740]*(10)+in_buf[741]*(18)+in_buf[742]*(48)+in_buf[743]*(3)+in_buf[744]*(6)+in_buf[745]*(51)+in_buf[746]*(48)+in_buf[747]*(39)+in_buf[748]*(68)+in_buf[749]*(49)+in_buf[750]*(29)+in_buf[751]*(1)+in_buf[752]*(10)+in_buf[753]*(-2)+in_buf[754]*(4)+in_buf[755]*(1)+in_buf[756]*(3)+in_buf[757]*(4)+in_buf[758]*(1)+in_buf[759]*(-3)+in_buf[760]*(-7)+in_buf[761]*(6)+in_buf[762]*(8)+in_buf[763]*(18)+in_buf[764]*(14)+in_buf[765]*(9)+in_buf[766]*(37)+in_buf[767]*(23)+in_buf[768]*(32)+in_buf[769]*(29)+in_buf[770]*(60)+in_buf[771]*(41)+in_buf[772]*(42)+in_buf[773]*(56)+in_buf[774]*(56)+in_buf[775]*(52)+in_buf[776]*(42)+in_buf[777]*(41)+in_buf[778]*(38)+in_buf[779]*(25)+in_buf[780]*(-1)+in_buf[781]*(4)+in_buf[782]*(-3)+in_buf[783]*(-3);
assign in_buf_weight049=in_buf[0]*(-3)+in_buf[1]*(-3)+in_buf[2]*(-3)+in_buf[3]*(2)+in_buf[4]*(0)+in_buf[5]*(-1)+in_buf[6]*(1)+in_buf[7]*(1)+in_buf[8]*(3)+in_buf[9]*(0)+in_buf[10]*(2)+in_buf[11]*(-2)+in_buf[12]*(-9)+in_buf[13]*(-4)+in_buf[14]*(21)+in_buf[15]*(11)+in_buf[16]*(2)+in_buf[17]*(-1)+in_buf[18]*(-3)+in_buf[19]*(2)+in_buf[20]*(3)+in_buf[21]*(3)+in_buf[22]*(3)+in_buf[23]*(0)+in_buf[24]*(3)+in_buf[25]*(3)+in_buf[26]*(-3)+in_buf[27]*(2)+in_buf[28]*(4)+in_buf[29]*(-3)+in_buf[30]*(0)+in_buf[31]*(1)+in_buf[32]*(-4)+in_buf[33]*(1)+in_buf[34]*(5)+in_buf[35]*(0)+in_buf[36]*(-4)+in_buf[37]*(-2)+in_buf[38]*(6)+in_buf[39]*(20)+in_buf[40]*(18)+in_buf[41]*(19)+in_buf[42]*(-12)+in_buf[43]*(7)+in_buf[44]*(41)+in_buf[45]*(26)+in_buf[46]*(-21)+in_buf[47]*(-21)+in_buf[48]*(-17)+in_buf[49]*(-15)+in_buf[50]*(-7)+in_buf[51]*(5)+in_buf[52]*(2)+in_buf[53]*(-3)+in_buf[54]*(1)+in_buf[55]*(-1)+in_buf[56]*(0)+in_buf[57]*(-2)+in_buf[58]*(-10)+in_buf[59]*(23)+in_buf[60]*(20)+in_buf[61]*(4)+in_buf[62]*(-4)+in_buf[63]*(9)+in_buf[64]*(24)+in_buf[65]*(39)+in_buf[66]*(61)+in_buf[67]*(37)+in_buf[68]*(8)+in_buf[69]*(-11)+in_buf[70]*(12)+in_buf[71]*(-10)+in_buf[72]*(-1)+in_buf[73]*(-17)+in_buf[74]*(-10)+in_buf[75]*(-17)+in_buf[76]*(2)+in_buf[77]*(25)+in_buf[78]*(18)+in_buf[79]*(14)+in_buf[80]*(14)+in_buf[81]*(16)+in_buf[82]*(3)+in_buf[83]*(-1)+in_buf[84]*(-1)+in_buf[85]*(-1)+in_buf[86]*(-13)+in_buf[87]*(27)+in_buf[88]*(-8)+in_buf[89]*(4)+in_buf[90]*(-5)+in_buf[91]*(-1)+in_buf[92]*(18)+in_buf[93]*(32)+in_buf[94]*(13)+in_buf[95]*(25)+in_buf[96]*(10)+in_buf[97]*(25)+in_buf[98]*(38)+in_buf[99]*(32)+in_buf[100]*(40)+in_buf[101]*(13)+in_buf[102]*(11)+in_buf[103]*(-13)+in_buf[104]*(-35)+in_buf[105]*(-3)+in_buf[106]*(-11)+in_buf[107]*(-2)+in_buf[108]*(-5)+in_buf[109]*(-15)+in_buf[110]*(-6)+in_buf[111]*(-2)+in_buf[112]*(-2)+in_buf[113]*(-1)+in_buf[114]*(-25)+in_buf[115]*(-26)+in_buf[116]*(-13)+in_buf[117]*(-3)+in_buf[118]*(1)+in_buf[119]*(15)+in_buf[120]*(13)+in_buf[121]*(12)+in_buf[122]*(-3)+in_buf[123]*(1)+in_buf[124]*(1)+in_buf[125]*(-12)+in_buf[126]*(0)+in_buf[127]*(14)+in_buf[128]*(38)+in_buf[129]*(31)+in_buf[130]*(3)+in_buf[131]*(9)+in_buf[132]*(9)+in_buf[133]*(-1)+in_buf[134]*(-7)+in_buf[135]*(-20)+in_buf[136]*(-9)+in_buf[137]*(10)+in_buf[138]*(10)+in_buf[139]*(30)+in_buf[140]*(-2)+in_buf[141]*(1)+in_buf[142]*(-29)+in_buf[143]*(8)+in_buf[144]*(14)+in_buf[145]*(-26)+in_buf[146]*(7)+in_buf[147]*(16)+in_buf[148]*(-8)+in_buf[149]*(-19)+in_buf[150]*(-16)+in_buf[151]*(-23)+in_buf[152]*(-13)+in_buf[153]*(-7)+in_buf[154]*(10)+in_buf[155]*(19)+in_buf[156]*(24)+in_buf[157]*(21)+in_buf[158]*(14)+in_buf[159]*(25)+in_buf[160]*(20)+in_buf[161]*(6)+in_buf[162]*(-10)+in_buf[163]*(-15)+in_buf[164]*(-15)+in_buf[165]*(-2)+in_buf[166]*(-11)+in_buf[167]*(15)+in_buf[168]*(-3)+in_buf[169]*(20)+in_buf[170]*(6)+in_buf[171]*(1)+in_buf[172]*(21)+in_buf[173]*(-13)+in_buf[174]*(6)+in_buf[175]*(7)+in_buf[176]*(-31)+in_buf[177]*(-33)+in_buf[178]*(-14)+in_buf[179]*(-21)+in_buf[180]*(-15)+in_buf[181]*(-5)+in_buf[182]*(4)+in_buf[183]*(6)+in_buf[184]*(7)+in_buf[185]*(-6)+in_buf[186]*(-11)+in_buf[187]*(2)+in_buf[188]*(-7)+in_buf[189]*(19)+in_buf[190]*(20)+in_buf[191]*(6)+in_buf[192]*(-19)+in_buf[193]*(-26)+in_buf[194]*(-27)+in_buf[195]*(-25)+in_buf[196]*(-2)+in_buf[197]*(23)+in_buf[198]*(4)+in_buf[199]*(-13)+in_buf[200]*(40)+in_buf[201]*(14)+in_buf[202]*(28)+in_buf[203]*(3)+in_buf[204]*(-14)+in_buf[205]*(-12)+in_buf[206]*(-9)+in_buf[207]*(12)+in_buf[208]*(0)+in_buf[209]*(9)+in_buf[210]*(-3)+in_buf[211]*(0)+in_buf[212]*(-14)+in_buf[213]*(-14)+in_buf[214]*(-1)+in_buf[215]*(-5)+in_buf[216]*(-12)+in_buf[217]*(13)+in_buf[218]*(30)+in_buf[219]*(8)+in_buf[220]*(3)+in_buf[221]*(23)+in_buf[222]*(-31)+in_buf[223]*(-39)+in_buf[224]*(31)+in_buf[225]*(4)+in_buf[226]*(-13)+in_buf[227]*(9)+in_buf[228]*(26)+in_buf[229]*(0)+in_buf[230]*(26)+in_buf[231]*(-4)+in_buf[232]*(-22)+in_buf[233]*(-6)+in_buf[234]*(7)+in_buf[235]*(12)+in_buf[236]*(19)+in_buf[237]*(24)+in_buf[238]*(22)+in_buf[239]*(13)+in_buf[240]*(2)+in_buf[241]*(-13)+in_buf[242]*(0)+in_buf[243]*(9)+in_buf[244]*(0)+in_buf[245]*(1)+in_buf[246]*(11)+in_buf[247]*(25)+in_buf[248]*(10)+in_buf[249]*(10)+in_buf[250]*(-4)+in_buf[251]*(1)+in_buf[252]*(3)+in_buf[253]*(-9)+in_buf[254]*(-28)+in_buf[255]*(23)+in_buf[256]*(26)+in_buf[257]*(18)+in_buf[258]*(12)+in_buf[259]*(-6)+in_buf[260]*(-20)+in_buf[261]*(-15)+in_buf[262]*(-11)+in_buf[263]*(-3)+in_buf[264]*(-1)+in_buf[265]*(22)+in_buf[266]*(14)+in_buf[267]*(-5)+in_buf[268]*(-20)+in_buf[269]*(-17)+in_buf[270]*(-7)+in_buf[271]*(9)+in_buf[272]*(13)+in_buf[273]*(4)+in_buf[274]*(-5)+in_buf[275]*(24)+in_buf[276]*(15)+in_buf[277]*(3)+in_buf[278]*(-22)+in_buf[279]*(-19)+in_buf[280]*(3)+in_buf[281]*(0)+in_buf[282]*(-5)+in_buf[283]*(19)+in_buf[284]*(17)+in_buf[285]*(27)+in_buf[286]*(30)+in_buf[287]*(1)+in_buf[288]*(-16)+in_buf[289]*(-21)+in_buf[290]*(-15)+in_buf[291]*(-4)+in_buf[292]*(-10)+in_buf[293]*(14)+in_buf[294]*(2)+in_buf[295]*(-28)+in_buf[296]*(-22)+in_buf[297]*(-1)+in_buf[298]*(5)+in_buf[299]*(-1)+in_buf[300]*(0)+in_buf[301]*(9)+in_buf[302]*(23)+in_buf[303]*(25)+in_buf[304]*(-6)+in_buf[305]*(-50)+in_buf[306]*(-4)+in_buf[307]*(-3)+in_buf[308]*(-9)+in_buf[309]*(23)+in_buf[310]*(1)+in_buf[311]*(17)+in_buf[312]*(8)+in_buf[313]*(3)+in_buf[314]*(17)+in_buf[315]*(18)+in_buf[316]*(-11)+in_buf[317]*(-8)+in_buf[318]*(-19)+in_buf[319]*(-14)+in_buf[320]*(7)+in_buf[321]*(7)+in_buf[322]*(3)+in_buf[323]*(-28)+in_buf[324]*(-31)+in_buf[325]*(-19)+in_buf[326]*(2)+in_buf[327]*(8)+in_buf[328]*(-7)+in_buf[329]*(12)+in_buf[330]*(14)+in_buf[331]*(10)+in_buf[332]*(-12)+in_buf[333]*(-3)+in_buf[334]*(12)+in_buf[335]*(-23)+in_buf[336]*(-14)+in_buf[337]*(0)+in_buf[338]*(10)+in_buf[339]*(8)+in_buf[340]*(6)+in_buf[341]*(-13)+in_buf[342]*(-11)+in_buf[343]*(-14)+in_buf[344]*(-25)+in_buf[345]*(-4)+in_buf[346]*(-29)+in_buf[347]*(-9)+in_buf[348]*(7)+in_buf[349]*(0)+in_buf[350]*(-8)+in_buf[351]*(-25)+in_buf[352]*(-27)+in_buf[353]*(-5)+in_buf[354]*(-15)+in_buf[355]*(0)+in_buf[356]*(1)+in_buf[357]*(11)+in_buf[358]*(13)+in_buf[359]*(7)+in_buf[360]*(28)+in_buf[361]*(20)+in_buf[362]*(3)+in_buf[363]*(-18)+in_buf[364]*(-1)+in_buf[365]*(13)+in_buf[366]*(22)+in_buf[367]*(5)+in_buf[368]*(-4)+in_buf[369]*(-19)+in_buf[370]*(-2)+in_buf[371]*(-16)+in_buf[372]*(-6)+in_buf[373]*(-12)+in_buf[374]*(-1)+in_buf[375]*(0)+in_buf[376]*(18)+in_buf[377]*(9)+in_buf[378]*(0)+in_buf[379]*(-13)+in_buf[380]*(-13)+in_buf[381]*(-11)+in_buf[382]*(-1)+in_buf[383]*(-4)+in_buf[384]*(-3)+in_buf[385]*(-9)+in_buf[386]*(18)+in_buf[387]*(25)+in_buf[388]*(38)+in_buf[389]*(61)+in_buf[390]*(59)+in_buf[391]*(28)+in_buf[392]*(0)+in_buf[393]*(9)+in_buf[394]*(19)+in_buf[395]*(-10)+in_buf[396]*(-3)+in_buf[397]*(4)+in_buf[398]*(2)+in_buf[399]*(3)+in_buf[400]*(-4)+in_buf[401]*(-11)+in_buf[402]*(0)+in_buf[403]*(13)+in_buf[404]*(13)+in_buf[405]*(5)+in_buf[406]*(-7)+in_buf[407]*(-2)+in_buf[408]*(-15)+in_buf[409]*(-14)+in_buf[410]*(-3)+in_buf[411]*(-5)+in_buf[412]*(-11)+in_buf[413]*(-3)+in_buf[414]*(18)+in_buf[415]*(6)+in_buf[416]*(27)+in_buf[417]*(58)+in_buf[418]*(53)+in_buf[419]*(17)+in_buf[420]*(1)+in_buf[421]*(-6)+in_buf[422]*(0)+in_buf[423]*(-4)+in_buf[424]*(0)+in_buf[425]*(0)+in_buf[426]*(0)+in_buf[427]*(12)+in_buf[428]*(10)+in_buf[429]*(6)+in_buf[430]*(9)+in_buf[431]*(14)+in_buf[432]*(8)+in_buf[433]*(4)+in_buf[434]*(3)+in_buf[435]*(-2)+in_buf[436]*(-4)+in_buf[437]*(-2)+in_buf[438]*(-2)+in_buf[439]*(2)+in_buf[440]*(1)+in_buf[441]*(0)+in_buf[442]*(18)+in_buf[443]*(2)+in_buf[444]*(32)+in_buf[445]*(39)+in_buf[446]*(14)+in_buf[447]*(44)+in_buf[448]*(0)+in_buf[449]*(-4)+in_buf[450]*(1)+in_buf[451]*(7)+in_buf[452]*(-2)+in_buf[453]*(1)+in_buf[454]*(7)+in_buf[455]*(24)+in_buf[456]*(35)+in_buf[457]*(26)+in_buf[458]*(31)+in_buf[459]*(23)+in_buf[460]*(8)+in_buf[461]*(-6)+in_buf[462]*(2)+in_buf[463]*(14)+in_buf[464]*(10)+in_buf[465]*(25)+in_buf[466]*(7)+in_buf[467]*(-1)+in_buf[468]*(3)+in_buf[469]*(16)+in_buf[470]*(33)+in_buf[471]*(24)+in_buf[472]*(6)+in_buf[473]*(36)+in_buf[474]*(57)+in_buf[475]*(46)+in_buf[476]*(-2)+in_buf[477]*(-15)+in_buf[478]*(26)+in_buf[479]*(0)+in_buf[480]*(21)+in_buf[481]*(11)+in_buf[482]*(17)+in_buf[483]*(24)+in_buf[484]*(33)+in_buf[485]*(34)+in_buf[486]*(17)+in_buf[487]*(21)+in_buf[488]*(10)+in_buf[489]*(-10)+in_buf[490]*(-1)+in_buf[491]*(9)+in_buf[492]*(18)+in_buf[493]*(21)+in_buf[494]*(-3)+in_buf[495]*(-5)+in_buf[496]*(-16)+in_buf[497]*(7)+in_buf[498]*(25)+in_buf[499]*(16)+in_buf[500]*(-1)+in_buf[501]*(13)+in_buf[502]*(19)+in_buf[503]*(59)+in_buf[504]*(-8)+in_buf[505]*(-18)+in_buf[506]*(12)+in_buf[507]*(0)+in_buf[508]*(16)+in_buf[509]*(7)+in_buf[510]*(19)+in_buf[511]*(33)+in_buf[512]*(31)+in_buf[513]*(24)+in_buf[514]*(13)+in_buf[515]*(14)+in_buf[516]*(6)+in_buf[517]*(-14)+in_buf[518]*(-7)+in_buf[519]*(18)+in_buf[520]*(35)+in_buf[521]*(14)+in_buf[522]*(-5)+in_buf[523]*(-12)+in_buf[524]*(-9)+in_buf[525]*(2)+in_buf[526]*(16)+in_buf[527]*(20)+in_buf[528]*(-2)+in_buf[529]*(17)+in_buf[530]*(3)+in_buf[531]*(25)+in_buf[532]*(-18)+in_buf[533]*(-10)+in_buf[534]*(24)+in_buf[535]*(12)+in_buf[536]*(35)+in_buf[537]*(27)+in_buf[538]*(10)+in_buf[539]*(20)+in_buf[540]*(20)+in_buf[541]*(15)+in_buf[542]*(21)+in_buf[543]*(13)+in_buf[544]*(-13)+in_buf[545]*(-17)+in_buf[546]*(3)+in_buf[547]*(16)+in_buf[548]*(22)+in_buf[549]*(14)+in_buf[550]*(-9)+in_buf[551]*(-13)+in_buf[552]*(-8)+in_buf[553]*(5)+in_buf[554]*(32)+in_buf[555]*(18)+in_buf[556]*(-13)+in_buf[557]*(5)+in_buf[558]*(63)+in_buf[559]*(8)+in_buf[560]*(1)+in_buf[561]*(22)+in_buf[562]*(44)+in_buf[563]*(47)+in_buf[564]*(37)+in_buf[565]*(24)+in_buf[566]*(9)+in_buf[567]*(31)+in_buf[568]*(23)+in_buf[569]*(8)+in_buf[570]*(18)+in_buf[571]*(16)+in_buf[572]*(-7)+in_buf[573]*(-15)+in_buf[574]*(-16)+in_buf[575]*(10)+in_buf[576]*(3)+in_buf[577]*(-1)+in_buf[578]*(-12)+in_buf[579]*(-17)+in_buf[580]*(1)+in_buf[581]*(16)+in_buf[582]*(20)+in_buf[583]*(19)+in_buf[584]*(-31)+in_buf[585]*(-10)+in_buf[586]*(50)+in_buf[587]*(-7)+in_buf[588]*(-8)+in_buf[589]*(15)+in_buf[590]*(33)+in_buf[591]*(39)+in_buf[592]*(31)+in_buf[593]*(9)+in_buf[594]*(18)+in_buf[595]*(25)+in_buf[596]*(12)+in_buf[597]*(16)+in_buf[598]*(9)+in_buf[599]*(15)+in_buf[600]*(0)+in_buf[601]*(-3)+in_buf[602]*(-15)+in_buf[603]*(-1)+in_buf[604]*(-7)+in_buf[605]*(-4)+in_buf[606]*(-11)+in_buf[607]*(-15)+in_buf[608]*(-4)+in_buf[609]*(2)+in_buf[610]*(54)+in_buf[611]*(22)+in_buf[612]*(-25)+in_buf[613]*(-16)+in_buf[614]*(37)+in_buf[615]*(6)+in_buf[616]*(-4)+in_buf[617]*(6)+in_buf[618]*(44)+in_buf[619]*(23)+in_buf[620]*(16)+in_buf[621]*(5)+in_buf[622]*(23)+in_buf[623]*(29)+in_buf[624]*(16)+in_buf[625]*(21)+in_buf[626]*(25)+in_buf[627]*(38)+in_buf[628]*(20)+in_buf[629]*(13)+in_buf[630]*(-8)+in_buf[631]*(-10)+in_buf[632]*(-15)+in_buf[633]*(-21)+in_buf[634]*(-18)+in_buf[635]*(0)+in_buf[636]*(-3)+in_buf[637]*(9)+in_buf[638]*(43)+in_buf[639]*(6)+in_buf[640]*(-9)+in_buf[641]*(-18)+in_buf[642]*(-19)+in_buf[643]*(0)+in_buf[644]*(-1)+in_buf[645]*(-3)+in_buf[646]*(36)+in_buf[647]*(35)+in_buf[648]*(11)+in_buf[649]*(-2)+in_buf[650]*(7)+in_buf[651]*(23)+in_buf[652]*(21)+in_buf[653]*(13)+in_buf[654]*(29)+in_buf[655]*(33)+in_buf[656]*(15)+in_buf[657]*(13)+in_buf[658]*(-1)+in_buf[659]*(-9)+in_buf[660]*(-22)+in_buf[661]*(-15)+in_buf[662]*(-1)+in_buf[663]*(-6)+in_buf[664]*(-20)+in_buf[665]*(-4)+in_buf[666]*(6)+in_buf[667]*(12)+in_buf[668]*(-22)+in_buf[669]*(-14)+in_buf[670]*(-37)+in_buf[671]*(0)+in_buf[672]*(-3)+in_buf[673]*(0)+in_buf[674]*(11)+in_buf[675]*(9)+in_buf[676]*(-3)+in_buf[677]*(-11)+in_buf[678]*(-12)+in_buf[679]*(-13)+in_buf[680]*(0)+in_buf[681]*(9)+in_buf[682]*(2)+in_buf[683]*(13)+in_buf[684]*(12)+in_buf[685]*(11)+in_buf[686]*(-2)+in_buf[687]*(0)+in_buf[688]*(3)+in_buf[689]*(-14)+in_buf[690]*(-8)+in_buf[691]*(-26)+in_buf[692]*(-24)+in_buf[693]*(-28)+in_buf[694]*(-17)+in_buf[695]*(-3)+in_buf[696]*(12)+in_buf[697]*(-1)+in_buf[698]*(-1)+in_buf[699]*(-2)+in_buf[700]*(4)+in_buf[701]*(2)+in_buf[702]*(-20)+in_buf[703]*(-17)+in_buf[704]*(-19)+in_buf[705]*(-55)+in_buf[706]*(-19)+in_buf[707]*(-13)+in_buf[708]*(-11)+in_buf[709]*(-11)+in_buf[710]*(22)+in_buf[711]*(-1)+in_buf[712]*(-42)+in_buf[713]*(-21)+in_buf[714]*(-4)+in_buf[715]*(-1)+in_buf[716]*(-2)+in_buf[717]*(-18)+in_buf[718]*(-35)+in_buf[719]*(-34)+in_buf[720]*(-41)+in_buf[721]*(-40)+in_buf[722]*(-34)+in_buf[723]*(-16)+in_buf[724]*(-21)+in_buf[725]*(3)+in_buf[726]*(16)+in_buf[727]*(4)+in_buf[728]*(3)+in_buf[729]*(4)+in_buf[730]*(-3)+in_buf[731]*(-3)+in_buf[732]*(-22)+in_buf[733]*(-48)+in_buf[734]*(-64)+in_buf[735]*(-41)+in_buf[736]*(2)+in_buf[737]*(-38)+in_buf[738]*(-41)+in_buf[739]*(-6)+in_buf[740]*(2)+in_buf[741]*(-9)+in_buf[742]*(-41)+in_buf[743]*(-54)+in_buf[744]*(-18)+in_buf[745]*(-32)+in_buf[746]*(-31)+in_buf[747]*(-24)+in_buf[748]*(-34)+in_buf[749]*(-25)+in_buf[750]*(-19)+in_buf[751]*(14)+in_buf[752]*(-14)+in_buf[753]*(5)+in_buf[754]*(2)+in_buf[755]*(3)+in_buf[756]*(-1)+in_buf[757]*(1)+in_buf[758]*(-3)+in_buf[759]*(4)+in_buf[760]*(1)+in_buf[761]*(2)+in_buf[762]*(0)+in_buf[763]*(2)+in_buf[764]*(-3)+in_buf[765]*(-17)+in_buf[766]*(-11)+in_buf[767]*(-20)+in_buf[768]*(-21)+in_buf[769]*(-11)+in_buf[770]*(-22)+in_buf[771]*(-12)+in_buf[772]*(-8)+in_buf[773]*(-30)+in_buf[774]*(-36)+in_buf[775]*(-4)+in_buf[776]*(-12)+in_buf[777]*(-29)+in_buf[778]*(-25)+in_buf[779]*(-21)+in_buf[780]*(3)+in_buf[781]*(2)+in_buf[782]*(-3)+in_buf[783]*(2);
assign in_buf_weight050=in_buf[0]*(3)+in_buf[1]*(-3)+in_buf[2]*(3)+in_buf[3]*(2)+in_buf[4]*(3)+in_buf[5]*(4)+in_buf[6]*(2)+in_buf[7]*(1)+in_buf[8]*(-3)+in_buf[9]*(2)+in_buf[10]*(-3)+in_buf[11]*(-2)+in_buf[12]*(7)+in_buf[13]*(9)+in_buf[14]*(-6)+in_buf[15]*(-3)+in_buf[16]*(-3)+in_buf[17]*(1)+in_buf[18]*(0)+in_buf[19]*(-1)+in_buf[20]*(3)+in_buf[21]*(0)+in_buf[22]*(-2)+in_buf[23]*(-2)+in_buf[24]*(-1)+in_buf[25]*(0)+in_buf[26]*(-3)+in_buf[27]*(-1)+in_buf[28]*(1)+in_buf[29]*(0)+in_buf[30]*(2)+in_buf[31]*(4)+in_buf[32]*(9)+in_buf[33]*(4)+in_buf[34]*(11)+in_buf[35]*(8)+in_buf[36]*(10)+in_buf[37]*(12)+in_buf[38]*(22)+in_buf[39]*(25)+in_buf[40]*(29)+in_buf[41]*(36)+in_buf[42]*(0)+in_buf[43]*(13)+in_buf[44]*(13)+in_buf[45]*(25)+in_buf[46]*(28)+in_buf[47]*(30)+in_buf[48]*(37)+in_buf[49]*(24)+in_buf[50]*(16)+in_buf[51]*(4)+in_buf[52]*(4)+in_buf[53]*(3)+in_buf[54]*(-1)+in_buf[55]*(1)+in_buf[56]*(-1)+in_buf[57]*(1)+in_buf[58]*(15)+in_buf[59]*(18)+in_buf[60]*(28)+in_buf[61]*(9)+in_buf[62]*(13)+in_buf[63]*(19)+in_buf[64]*(5)+in_buf[65]*(-16)+in_buf[66]*(-11)+in_buf[67]*(14)+in_buf[68]*(2)+in_buf[69]*(-12)+in_buf[70]*(-14)+in_buf[71]*(2)+in_buf[72]*(19)+in_buf[73]*(16)+in_buf[74]*(26)+in_buf[75]*(19)+in_buf[76]*(12)+in_buf[77]*(19)+in_buf[78]*(35)+in_buf[79]*(16)+in_buf[80]*(-8)+in_buf[81]*(-10)+in_buf[82]*(2)+in_buf[83]*(-2)+in_buf[84]*(2)+in_buf[85]*(-2)+in_buf[86]*(-15)+in_buf[87]*(26)+in_buf[88]*(31)+in_buf[89]*(-4)+in_buf[90]*(0)+in_buf[91]*(3)+in_buf[92]*(-12)+in_buf[93]*(-12)+in_buf[94]*(-25)+in_buf[95]*(3)+in_buf[96]*(5)+in_buf[97]*(8)+in_buf[98]*(4)+in_buf[99]*(-2)+in_buf[100]*(-5)+in_buf[101]*(8)+in_buf[102]*(15)+in_buf[103]*(17)+in_buf[104]*(6)+in_buf[105]*(18)+in_buf[106]*(21)+in_buf[107]*(26)+in_buf[108]*(15)+in_buf[109]*(-19)+in_buf[110]*(7)+in_buf[111]*(0)+in_buf[112]*(1)+in_buf[113]*(-2)+in_buf[114]*(-17)+in_buf[115]*(-5)+in_buf[116]*(-18)+in_buf[117]*(-30)+in_buf[118]*(-24)+in_buf[119]*(-24)+in_buf[120]*(-34)+in_buf[121]*(-36)+in_buf[122]*(-15)+in_buf[123]*(-13)+in_buf[124]*(-10)+in_buf[125]*(-11)+in_buf[126]*(-16)+in_buf[127]*(-14)+in_buf[128]*(-13)+in_buf[129]*(1)+in_buf[130]*(-3)+in_buf[131]*(8)+in_buf[132]*(5)+in_buf[133]*(12)+in_buf[134]*(-6)+in_buf[135]*(25)+in_buf[136]*(16)+in_buf[137]*(24)+in_buf[138]*(20)+in_buf[139]*(24)+in_buf[140]*(-2)+in_buf[141]*(1)+in_buf[142]*(20)+in_buf[143]*(-10)+in_buf[144]*(-23)+in_buf[145]*(-33)+in_buf[146]*(-38)+in_buf[147]*(-32)+in_buf[148]*(-25)+in_buf[149]*(6)+in_buf[150]*(13)+in_buf[151]*(0)+in_buf[152]*(-1)+in_buf[153]*(-5)+in_buf[154]*(2)+in_buf[155]*(-7)+in_buf[156]*(1)+in_buf[157]*(11)+in_buf[158]*(-5)+in_buf[159]*(-8)+in_buf[160]*(5)+in_buf[161]*(9)+in_buf[162]*(-1)+in_buf[163]*(10)+in_buf[164]*(21)+in_buf[165]*(27)+in_buf[166]*(44)+in_buf[167]*(19)+in_buf[168]*(-3)+in_buf[169]*(20)+in_buf[170]*(29)+in_buf[171]*(-27)+in_buf[172]*(-18)+in_buf[173]*(-14)+in_buf[174]*(-57)+in_buf[175]*(-23)+in_buf[176]*(-10)+in_buf[177]*(-12)+in_buf[178]*(1)+in_buf[179]*(0)+in_buf[180]*(-1)+in_buf[181]*(-2)+in_buf[182]*(0)+in_buf[183]*(-4)+in_buf[184]*(-6)+in_buf[185]*(-4)+in_buf[186]*(-11)+in_buf[187]*(-7)+in_buf[188]*(-25)+in_buf[189]*(-21)+in_buf[190]*(17)+in_buf[191]*(7)+in_buf[192]*(32)+in_buf[193]*(51)+in_buf[194]*(21)+in_buf[195]*(26)+in_buf[196]*(-1)+in_buf[197]*(-3)+in_buf[198]*(25)+in_buf[199]*(-28)+in_buf[200]*(-32)+in_buf[201]*(-34)+in_buf[202]*(-54)+in_buf[203]*(-48)+in_buf[204]*(-12)+in_buf[205]*(10)+in_buf[206]*(3)+in_buf[207]*(6)+in_buf[208]*(0)+in_buf[209]*(-2)+in_buf[210]*(-6)+in_buf[211]*(-5)+in_buf[212]*(-7)+in_buf[213]*(-7)+in_buf[214]*(0)+in_buf[215]*(-10)+in_buf[216]*(-19)+in_buf[217]*(-13)+in_buf[218]*(12)+in_buf[219]*(14)+in_buf[220]*(17)+in_buf[221]*(27)+in_buf[222]*(35)+in_buf[223]*(35)+in_buf[224]*(14)+in_buf[225]*(-27)+in_buf[226]*(20)+in_buf[227]*(-15)+in_buf[228]*(-35)+in_buf[229]*(-49)+in_buf[230]*(-38)+in_buf[231]*(-33)+in_buf[232]*(-14)+in_buf[233]*(18)+in_buf[234]*(0)+in_buf[235]*(10)+in_buf[236]*(7)+in_buf[237]*(1)+in_buf[238]*(-5)+in_buf[239]*(-13)+in_buf[240]*(-10)+in_buf[241]*(-8)+in_buf[242]*(-6)+in_buf[243]*(3)+in_buf[244]*(2)+in_buf[245]*(12)+in_buf[246]*(-1)+in_buf[247]*(7)+in_buf[248]*(22)+in_buf[249]*(16)+in_buf[250]*(-1)+in_buf[251]*(8)+in_buf[252]*(-5)+in_buf[253]*(-11)+in_buf[254]*(-4)+in_buf[255]*(-27)+in_buf[256]*(-38)+in_buf[257]*(-43)+in_buf[258]*(-24)+in_buf[259]*(-24)+in_buf[260]*(-10)+in_buf[261]*(8)+in_buf[262]*(4)+in_buf[263]*(12)+in_buf[264]*(0)+in_buf[265]*(0)+in_buf[266]*(-14)+in_buf[267]*(-32)+in_buf[268]*(-15)+in_buf[269]*(-10)+in_buf[270]*(-1)+in_buf[271]*(0)+in_buf[272]*(0)+in_buf[273]*(-6)+in_buf[274]*(-17)+in_buf[275]*(5)+in_buf[276]*(45)+in_buf[277]*(34)+in_buf[278]*(-8)+in_buf[279]*(-26)+in_buf[280]*(-7)+in_buf[281]*(-7)+in_buf[282]*(16)+in_buf[283]*(2)+in_buf[284]*(-2)+in_buf[285]*(-7)+in_buf[286]*(-19)+in_buf[287]*(-13)+in_buf[288]*(2)+in_buf[289]*(27)+in_buf[290]*(12)+in_buf[291]*(-2)+in_buf[292]*(3)+in_buf[293]*(3)+in_buf[294]*(-9)+in_buf[295]*(-11)+in_buf[296]*(-8)+in_buf[297]*(3)+in_buf[298]*(4)+in_buf[299]*(-3)+in_buf[300]*(-11)+in_buf[301]*(-11)+in_buf[302]*(-11)+in_buf[303]*(0)+in_buf[304]*(25)+in_buf[305]*(7)+in_buf[306]*(10)+in_buf[307]*(-34)+in_buf[308]*(0)+in_buf[309]*(-3)+in_buf[310]*(11)+in_buf[311]*(-14)+in_buf[312]*(-9)+in_buf[313]*(-33)+in_buf[314]*(-19)+in_buf[315]*(-18)+in_buf[316]*(-1)+in_buf[317]*(12)+in_buf[318]*(8)+in_buf[319]*(1)+in_buf[320]*(0)+in_buf[321]*(-3)+in_buf[322]*(-7)+in_buf[323]*(-12)+in_buf[324]*(-8)+in_buf[325]*(-6)+in_buf[326]*(-1)+in_buf[327]*(-8)+in_buf[328]*(-35)+in_buf[329]*(-27)+in_buf[330]*(-30)+in_buf[331]*(-24)+in_buf[332]*(-14)+in_buf[333]*(0)+in_buf[334]*(27)+in_buf[335]*(-23)+in_buf[336]*(0)+in_buf[337]*(-1)+in_buf[338]*(8)+in_buf[339]*(-4)+in_buf[340]*(-26)+in_buf[341]*(-36)+in_buf[342]*(-34)+in_buf[343]*(-16)+in_buf[344]*(0)+in_buf[345]*(11)+in_buf[346]*(17)+in_buf[347]*(19)+in_buf[348]*(14)+in_buf[349]*(10)+in_buf[350]*(-9)+in_buf[351]*(-4)+in_buf[352]*(-12)+in_buf[353]*(-14)+in_buf[354]*(-7)+in_buf[355]*(-5)+in_buf[356]*(-13)+in_buf[357]*(-7)+in_buf[358]*(-19)+in_buf[359]*(-29)+in_buf[360]*(-12)+in_buf[361]*(0)+in_buf[362]*(24)+in_buf[363]*(-30)+in_buf[364]*(-1)+in_buf[365]*(-3)+in_buf[366]*(-7)+in_buf[367]*(-3)+in_buf[368]*(-38)+in_buf[369]*(-25)+in_buf[370]*(-17)+in_buf[371]*(2)+in_buf[372]*(-3)+in_buf[373]*(14)+in_buf[374]*(26)+in_buf[375]*(25)+in_buf[376]*(28)+in_buf[377]*(1)+in_buf[378]*(-6)+in_buf[379]*(4)+in_buf[380]*(-11)+in_buf[381]*(-6)+in_buf[382]*(2)+in_buf[383]*(7)+in_buf[384]*(1)+in_buf[385]*(9)+in_buf[386]*(4)+in_buf[387]*(5)+in_buf[388]*(-22)+in_buf[389]*(-15)+in_buf[390]*(-2)+in_buf[391]*(-2)+in_buf[392]*(17)+in_buf[393]*(-6)+in_buf[394]*(-4)+in_buf[395]*(-6)+in_buf[396]*(-39)+in_buf[397]*(-8)+in_buf[398]*(-11)+in_buf[399]*(-9)+in_buf[400]*(0)+in_buf[401]*(6)+in_buf[402]*(18)+in_buf[403]*(21)+in_buf[404]*(14)+in_buf[405]*(2)+in_buf[406]*(-3)+in_buf[407]*(-3)+in_buf[408]*(-20)+in_buf[409]*(-1)+in_buf[410]*(3)+in_buf[411]*(-10)+in_buf[412]*(19)+in_buf[413]*(32)+in_buf[414]*(5)+in_buf[415]*(-2)+in_buf[416]*(1)+in_buf[417]*(-2)+in_buf[418]*(-14)+in_buf[419]*(-14)+in_buf[420]*(13)+in_buf[421]*(1)+in_buf[422]*(3)+in_buf[423]*(-5)+in_buf[424]*(-26)+in_buf[425]*(-26)+in_buf[426]*(-15)+in_buf[427]*(-1)+in_buf[428]*(-5)+in_buf[429]*(13)+in_buf[430]*(9)+in_buf[431]*(18)+in_buf[432]*(19)+in_buf[433]*(-9)+in_buf[434]*(-1)+in_buf[435]*(-8)+in_buf[436]*(-16)+in_buf[437]*(2)+in_buf[438]*(0)+in_buf[439]*(-7)+in_buf[440]*(15)+in_buf[441]*(28)+in_buf[442]*(0)+in_buf[443]*(20)+in_buf[444]*(6)+in_buf[445]*(30)+in_buf[446]*(-19)+in_buf[447]*(-12)+in_buf[448]*(-5)+in_buf[449]*(0)+in_buf[450]*(-19)+in_buf[451]*(9)+in_buf[452]*(-23)+in_buf[453]*(-21)+in_buf[454]*(-13)+in_buf[455]*(1)+in_buf[456]*(5)+in_buf[457]*(5)+in_buf[458]*(7)+in_buf[459]*(14)+in_buf[460]*(11)+in_buf[461]*(1)+in_buf[462]*(6)+in_buf[463]*(0)+in_buf[464]*(-23)+in_buf[465]*(-3)+in_buf[466]*(3)+in_buf[467]*(11)+in_buf[468]*(12)+in_buf[469]*(21)+in_buf[470]*(24)+in_buf[471]*(3)+in_buf[472]*(-4)+in_buf[473]*(25)+in_buf[474]*(-29)+in_buf[475]*(-30)+in_buf[476]*(4)+in_buf[477]*(-3)+in_buf[478]*(-31)+in_buf[479]*(9)+in_buf[480]*(-4)+in_buf[481]*(1)+in_buf[482]*(0)+in_buf[483]*(-1)+in_buf[484]*(-1)+in_buf[485]*(0)+in_buf[486]*(0)+in_buf[487]*(0)+in_buf[488]*(0)+in_buf[489]*(-11)+in_buf[490]*(-10)+in_buf[491]*(4)+in_buf[492]*(-5)+in_buf[493]*(-1)+in_buf[494]*(3)+in_buf[495]*(10)+in_buf[496]*(3)+in_buf[497]*(12)+in_buf[498]*(5)+in_buf[499]*(-6)+in_buf[500]*(-34)+in_buf[501]*(-31)+in_buf[502]*(-56)+in_buf[503]*(1)+in_buf[504]*(-37)+in_buf[505]*(-13)+in_buf[506]*(-38)+in_buf[507]*(25)+in_buf[508]*(13)+in_buf[509]*(10)+in_buf[510]*(19)+in_buf[511]*(6)+in_buf[512]*(7)+in_buf[513]*(4)+in_buf[514]*(-5)+in_buf[515]*(-5)+in_buf[516]*(3)+in_buf[517]*(-15)+in_buf[518]*(-6)+in_buf[519]*(9)+in_buf[520]*(5)+in_buf[521]*(-10)+in_buf[522]*(-1)+in_buf[523]*(-1)+in_buf[524]*(-13)+in_buf[525]*(-4)+in_buf[526]*(-9)+in_buf[527]*(-21)+in_buf[528]*(-29)+in_buf[529]*(-24)+in_buf[530]*(-44)+in_buf[531]*(0)+in_buf[532]*(-3)+in_buf[533]*(-22)+in_buf[534]*(-18)+in_buf[535]*(19)+in_buf[536]*(11)+in_buf[537]*(-1)+in_buf[538]*(5)+in_buf[539]*(-1)+in_buf[540]*(11)+in_buf[541]*(14)+in_buf[542]*(15)+in_buf[543]*(17)+in_buf[544]*(-1)+in_buf[545]*(-19)+in_buf[546]*(0)+in_buf[547]*(15)+in_buf[548]*(8)+in_buf[549]*(2)+in_buf[550]*(5)+in_buf[551]*(-2)+in_buf[552]*(-1)+in_buf[553]*(0)+in_buf[554]*(2)+in_buf[555]*(-2)+in_buf[556]*(-12)+in_buf[557]*(-20)+in_buf[558]*(-7)+in_buf[559]*(5)+in_buf[560]*(0)+in_buf[561]*(22)+in_buf[562]*(-11)+in_buf[563]*(0)+in_buf[564]*(4)+in_buf[565]*(-6)+in_buf[566]*(-16)+in_buf[567]*(-3)+in_buf[568]*(22)+in_buf[569]*(35)+in_buf[570]*(32)+in_buf[571]*(23)+in_buf[572]*(3)+in_buf[573]*(1)+in_buf[574]*(0)+in_buf[575]*(11)+in_buf[576]*(-12)+in_buf[577]*(-6)+in_buf[578]*(-5)+in_buf[579]*(-7)+in_buf[580]*(0)+in_buf[581]*(1)+in_buf[582]*(15)+in_buf[583]*(-20)+in_buf[584]*(-22)+in_buf[585]*(-7)+in_buf[586]*(-16)+in_buf[587]*(0)+in_buf[588]*(-5)+in_buf[589]*(-9)+in_buf[590]*(-18)+in_buf[591]*(5)+in_buf[592]*(-8)+in_buf[593]*(-16)+in_buf[594]*(-27)+in_buf[595]*(-2)+in_buf[596]*(7)+in_buf[597]*(29)+in_buf[598]*(18)+in_buf[599]*(29)+in_buf[600]*(13)+in_buf[601]*(16)+in_buf[602]*(19)+in_buf[603]*(10)+in_buf[604]*(-5)+in_buf[605]*(6)+in_buf[606]*(-7)+in_buf[607]*(-8)+in_buf[608]*(-3)+in_buf[609]*(4)+in_buf[610]*(8)+in_buf[611]*(-22)+in_buf[612]*(-24)+in_buf[613]*(2)+in_buf[614]*(18)+in_buf[615]*(2)+in_buf[616]*(-8)+in_buf[617]*(-9)+in_buf[618]*(7)+in_buf[619]*(20)+in_buf[620]*(-15)+in_buf[621]*(-33)+in_buf[622]*(-29)+in_buf[623]*(-16)+in_buf[624]*(-10)+in_buf[625]*(13)+in_buf[626]*(27)+in_buf[627]*(40)+in_buf[628]*(26)+in_buf[629]*(14)+in_buf[630]*(-4)+in_buf[631]*(10)+in_buf[632]*(8)+in_buf[633]*(-7)+in_buf[634]*(-15)+in_buf[635]*(-4)+in_buf[636]*(-8)+in_buf[637]*(-2)+in_buf[638]*(0)+in_buf[639]*(-7)+in_buf[640]*(-7)+in_buf[641]*(-2)+in_buf[642]*(18)+in_buf[643]*(-5)+in_buf[644]*(-2)+in_buf[645]*(1)+in_buf[646]*(12)+in_buf[647]*(35)+in_buf[648]*(16)+in_buf[649]*(-20)+in_buf[650]*(-4)+in_buf[651]*(-5)+in_buf[652]*(16)+in_buf[653]*(11)+in_buf[654]*(18)+in_buf[655]*(17)+in_buf[656]*(16)+in_buf[657]*(6)+in_buf[658]*(2)+in_buf[659]*(-1)+in_buf[660]*(0)+in_buf[661]*(-16)+in_buf[662]*(-20)+in_buf[663]*(-25)+in_buf[664]*(-22)+in_buf[665]*(-15)+in_buf[666]*(-16)+in_buf[667]*(2)+in_buf[668]*(-9)+in_buf[669]*(4)+in_buf[670]*(0)+in_buf[671]*(4)+in_buf[672]*(3)+in_buf[673]*(-2)+in_buf[674]*(-10)+in_buf[675]*(6)+in_buf[676]*(-5)+in_buf[677]*(-11)+in_buf[678]*(-7)+in_buf[679]*(-9)+in_buf[680]*(-1)+in_buf[681]*(7)+in_buf[682]*(-1)+in_buf[683]*(3)+in_buf[684]*(6)+in_buf[685]*(12)+in_buf[686]*(23)+in_buf[687]*(12)+in_buf[688]*(13)+in_buf[689]*(-14)+in_buf[690]*(-24)+in_buf[691]*(-38)+in_buf[692]*(-27)+in_buf[693]*(-27)+in_buf[694]*(-6)+in_buf[695]*(-8)+in_buf[696]*(0)+in_buf[697]*(-21)+in_buf[698]*(-17)+in_buf[699]*(-1)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(4)+in_buf[703]*(8)+in_buf[704]*(-16)+in_buf[705]*(-34)+in_buf[706]*(-15)+in_buf[707]*(-18)+in_buf[708]*(-46)+in_buf[709]*(-34)+in_buf[710]*(-3)+in_buf[711]*(0)+in_buf[712]*(-19)+in_buf[713]*(0)+in_buf[714]*(-4)+in_buf[715]*(13)+in_buf[716]*(-6)+in_buf[717]*(-31)+in_buf[718]*(-21)+in_buf[719]*(7)+in_buf[720]*(-11)+in_buf[721]*(-7)+in_buf[722]*(3)+in_buf[723]*(19)+in_buf[724]*(13)+in_buf[725]*(1)+in_buf[726]*(1)+in_buf[727]*(-1)+in_buf[728]*(0)+in_buf[729]*(4)+in_buf[730]*(-2)+in_buf[731]*(-1)+in_buf[732]*(-13)+in_buf[733]*(-22)+in_buf[734]*(-45)+in_buf[735]*(-41)+in_buf[736]*(-43)+in_buf[737]*(-53)+in_buf[738]*(-36)+in_buf[739]*(9)+in_buf[740]*(8)+in_buf[741]*(15)+in_buf[742]*(-23)+in_buf[743]*(-18)+in_buf[744]*(-17)+in_buf[745]*(-19)+in_buf[746]*(-10)+in_buf[747]*(8)+in_buf[748]*(8)+in_buf[749]*(8)+in_buf[750]*(9)+in_buf[751]*(21)+in_buf[752]*(9)+in_buf[753]*(0)+in_buf[754]*(1)+in_buf[755]*(0)+in_buf[756]*(2)+in_buf[757]*(2)+in_buf[758]*(3)+in_buf[759]*(2)+in_buf[760]*(-5)+in_buf[761]*(-2)+in_buf[762]*(-4)+in_buf[763]*(-3)+in_buf[764]*(-5)+in_buf[765]*(-2)+in_buf[766]*(-25)+in_buf[767]*(-13)+in_buf[768]*(-1)+in_buf[769]*(0)+in_buf[770]*(-19)+in_buf[771]*(-13)+in_buf[772]*(-6)+in_buf[773]*(-5)+in_buf[774]*(0)+in_buf[775]*(-17)+in_buf[776]*(-12)+in_buf[777]*(-20)+in_buf[778]*(-13)+in_buf[779]*(-5)+in_buf[780]*(-2)+in_buf[781]*(-3)+in_buf[782]*(-3)+in_buf[783]*(3);
assign in_buf_weight051=in_buf[0]*(2)+in_buf[1]*(4)+in_buf[2]*(0)+in_buf[3]*(-2)+in_buf[4]*(0)+in_buf[5]*(2)+in_buf[6]*(-1)+in_buf[7]*(-1)+in_buf[8]*(1)+in_buf[9]*(4)+in_buf[10]*(-3)+in_buf[11]*(0)+in_buf[12]*(10)+in_buf[13]*(8)+in_buf[14]*(-16)+in_buf[15]*(-18)+in_buf[16]*(-3)+in_buf[17]*(1)+in_buf[18]*(0)+in_buf[19]*(4)+in_buf[20]*(-3)+in_buf[21]*(1)+in_buf[22]*(0)+in_buf[23]*(4)+in_buf[24]*(0)+in_buf[25]*(4)+in_buf[26]*(4)+in_buf[27]*(1)+in_buf[28]*(0)+in_buf[29]*(0)+in_buf[30]*(1)+in_buf[31]*(0)+in_buf[32]*(9)+in_buf[33]*(0)+in_buf[34]*(-1)+in_buf[35]*(-1)+in_buf[36]*(6)+in_buf[37]*(11)+in_buf[38]*(23)+in_buf[39]*(-6)+in_buf[40]*(-10)+in_buf[41]*(-2)+in_buf[42]*(7)+in_buf[43]*(-26)+in_buf[44]*(-32)+in_buf[45]*(-23)+in_buf[46]*(31)+in_buf[47]*(24)+in_buf[48]*(37)+in_buf[49]*(31)+in_buf[50]*(21)+in_buf[51]*(12)+in_buf[52]*(0)+in_buf[53]*(1)+in_buf[54]*(-3)+in_buf[55]*(3)+in_buf[56]*(0)+in_buf[57]*(5)+in_buf[58]*(5)+in_buf[59]*(-4)+in_buf[60]*(8)+in_buf[61]*(0)+in_buf[62]*(12)+in_buf[63]*(9)+in_buf[64]*(3)+in_buf[65]*(-17)+in_buf[66]*(-16)+in_buf[67]*(5)+in_buf[68]*(-1)+in_buf[69]*(-9)+in_buf[70]*(-26)+in_buf[71]*(-8)+in_buf[72]*(-1)+in_buf[73]*(17)+in_buf[74]*(16)+in_buf[75]*(26)+in_buf[76]*(16)+in_buf[77]*(18)+in_buf[78]*(13)+in_buf[79]*(-5)+in_buf[80]*(9)+in_buf[81]*(2)+in_buf[82]*(-3)+in_buf[83]*(0)+in_buf[84]*(2)+in_buf[85]*(0)+in_buf[86]*(-6)+in_buf[87]*(-2)+in_buf[88]*(2)+in_buf[89]*(2)+in_buf[90]*(11)+in_buf[91]*(21)+in_buf[92]*(-2)+in_buf[93]*(-49)+in_buf[94]*(-17)+in_buf[95]*(-15)+in_buf[96]*(-26)+in_buf[97]*(-23)+in_buf[98]*(-19)+in_buf[99]*(3)+in_buf[100]*(1)+in_buf[101]*(1)+in_buf[102]*(-2)+in_buf[103]*(6)+in_buf[104]*(8)+in_buf[105]*(22)+in_buf[106]*(24)+in_buf[107]*(28)+in_buf[108]*(-3)+in_buf[109]*(-18)+in_buf[110]*(-11)+in_buf[111]*(3)+in_buf[112]*(-2)+in_buf[113]*(4)+in_buf[114]*(6)+in_buf[115]*(24)+in_buf[116]*(46)+in_buf[117]*(33)+in_buf[118]*(6)+in_buf[119]*(10)+in_buf[120]*(29)+in_buf[121]*(3)+in_buf[122]*(-2)+in_buf[123]*(-15)+in_buf[124]*(-17)+in_buf[125]*(3)+in_buf[126]*(-2)+in_buf[127]*(-4)+in_buf[128]*(5)+in_buf[129]*(0)+in_buf[130]*(-12)+in_buf[131]*(1)+in_buf[132]*(0)+in_buf[133]*(0)+in_buf[134]*(28)+in_buf[135]*(13)+in_buf[136]*(10)+in_buf[137]*(-22)+in_buf[138]*(-33)+in_buf[139]*(16)+in_buf[140]*(-1)+in_buf[141]*(-1)+in_buf[142]*(8)+in_buf[143]*(16)+in_buf[144]*(20)+in_buf[145]*(38)+in_buf[146]*(25)+in_buf[147]*(20)+in_buf[148]*(-2)+in_buf[149]*(-13)+in_buf[150]*(-29)+in_buf[151]*(-28)+in_buf[152]*(-2)+in_buf[153]*(6)+in_buf[154]*(4)+in_buf[155]*(5)+in_buf[156]*(-13)+in_buf[157]*(-9)+in_buf[158]*(0)+in_buf[159]*(16)+in_buf[160]*(-3)+in_buf[161]*(1)+in_buf[162]*(0)+in_buf[163]*(26)+in_buf[164]*(34)+in_buf[165]*(18)+in_buf[166]*(-9)+in_buf[167]*(17)+in_buf[168]*(1)+in_buf[169]*(26)+in_buf[170]*(1)+in_buf[171]*(-1)+in_buf[172]*(-10)+in_buf[173]*(0)+in_buf[174]*(13)+in_buf[175]*(4)+in_buf[176]*(-4)+in_buf[177]*(-2)+in_buf[178]*(-3)+in_buf[179]*(-4)+in_buf[180]*(-1)+in_buf[181]*(9)+in_buf[182]*(2)+in_buf[183]*(-2)+in_buf[184]*(-6)+in_buf[185]*(-10)+in_buf[186]*(-14)+in_buf[187]*(-12)+in_buf[188]*(9)+in_buf[189]*(16)+in_buf[190]*(-9)+in_buf[191]*(8)+in_buf[192]*(1)+in_buf[193]*(14)+in_buf[194]*(6)+in_buf[195]*(6)+in_buf[196]*(4)+in_buf[197]*(18)+in_buf[198]*(-14)+in_buf[199]*(-11)+in_buf[200]*(22)+in_buf[201]*(1)+in_buf[202]*(5)+in_buf[203]*(-6)+in_buf[204]*(-7)+in_buf[205]*(0)+in_buf[206]*(2)+in_buf[207]*(-10)+in_buf[208]*(0)+in_buf[209]*(-3)+in_buf[210]*(-1)+in_buf[211]*(-1)+in_buf[212]*(-7)+in_buf[213]*(-9)+in_buf[214]*(-12)+in_buf[215]*(-10)+in_buf[216]*(1)+in_buf[217]*(0)+in_buf[218]*(-6)+in_buf[219]*(-10)+in_buf[220]*(-17)+in_buf[221]*(1)+in_buf[222]*(-20)+in_buf[223]*(-3)+in_buf[224]*(-4)+in_buf[225]*(-29)+in_buf[226]*(14)+in_buf[227]*(33)+in_buf[228]*(20)+in_buf[229]*(26)+in_buf[230]*(5)+in_buf[231]*(-10)+in_buf[232]*(-7)+in_buf[233]*(-10)+in_buf[234]*(-12)+in_buf[235]*(-20)+in_buf[236]*(-18)+in_buf[237]*(-3)+in_buf[238]*(-9)+in_buf[239]*(-1)+in_buf[240]*(-3)+in_buf[241]*(0)+in_buf[242]*(2)+in_buf[243]*(0)+in_buf[244]*(-3)+in_buf[245]*(9)+in_buf[246]*(-8)+in_buf[247]*(-30)+in_buf[248]*(-58)+in_buf[249]*(-42)+in_buf[250]*(-17)+in_buf[251]*(-18)+in_buf[252]*(-6)+in_buf[253]*(-27)+in_buf[254]*(17)+in_buf[255]*(4)+in_buf[256]*(16)+in_buf[257]*(19)+in_buf[258]*(3)+in_buf[259]*(1)+in_buf[260]*(3)+in_buf[261]*(4)+in_buf[262]*(-17)+in_buf[263]*(-27)+in_buf[264]*(-18)+in_buf[265]*(-4)+in_buf[266]*(3)+in_buf[267]*(5)+in_buf[268]*(9)+in_buf[269]*(14)+in_buf[270]*(13)+in_buf[271]*(13)+in_buf[272]*(9)+in_buf[273]*(-2)+in_buf[274]*(-37)+in_buf[275]*(-48)+in_buf[276]*(-62)+in_buf[277]*(-52)+in_buf[278]*(-42)+in_buf[279]*(-33)+in_buf[280]*(-8)+in_buf[281]*(-14)+in_buf[282]*(-16)+in_buf[283]*(8)+in_buf[284]*(0)+in_buf[285]*(10)+in_buf[286]*(-3)+in_buf[287]*(0)+in_buf[288]*(0)+in_buf[289]*(-11)+in_buf[290]*(-23)+in_buf[291]*(-20)+in_buf[292]*(-7)+in_buf[293]*(6)+in_buf[294]*(1)+in_buf[295]*(-4)+in_buf[296]*(6)+in_buf[297]*(20)+in_buf[298]*(22)+in_buf[299]*(20)+in_buf[300]*(-3)+in_buf[301]*(-20)+in_buf[302]*(-51)+in_buf[303]*(-45)+in_buf[304]*(-75)+in_buf[305]*(-50)+in_buf[306]*(-27)+in_buf[307]*(-10)+in_buf[308]*(-1)+in_buf[309]*(-24)+in_buf[310]*(-19)+in_buf[311]*(22)+in_buf[312]*(4)+in_buf[313]*(15)+in_buf[314]*(-11)+in_buf[315]*(-4)+in_buf[316]*(-1)+in_buf[317]*(-7)+in_buf[318]*(-5)+in_buf[319]*(0)+in_buf[320]*(20)+in_buf[321]*(20)+in_buf[322]*(22)+in_buf[323]*(13)+in_buf[324]*(3)+in_buf[325]*(11)+in_buf[326]*(14)+in_buf[327]*(10)+in_buf[328]*(5)+in_buf[329]*(-17)+in_buf[330]*(-41)+in_buf[331]*(-56)+in_buf[332]*(-76)+in_buf[333]*(-69)+in_buf[334]*(-33)+in_buf[335]*(-13)+in_buf[336]*(0)+in_buf[337]*(2)+in_buf[338]*(-19)+in_buf[339]*(-6)+in_buf[340]*(10)+in_buf[341]*(25)+in_buf[342]*(1)+in_buf[343]*(-4)+in_buf[344]*(-17)+in_buf[345]*(-4)+in_buf[346]*(6)+in_buf[347]*(19)+in_buf[348]*(30)+in_buf[349]*(36)+in_buf[350]*(24)+in_buf[351]*(14)+in_buf[352]*(18)+in_buf[353]*(14)+in_buf[354]*(11)+in_buf[355]*(5)+in_buf[356]*(-6)+in_buf[357]*(-12)+in_buf[358]*(-26)+in_buf[359]*(-8)+in_buf[360]*(-19)+in_buf[361]*(-59)+in_buf[362]*(-52)+in_buf[363]*(-34)+in_buf[364]*(16)+in_buf[365]*(0)+in_buf[366]*(-19)+in_buf[367]*(-8)+in_buf[368]*(14)+in_buf[369]*(3)+in_buf[370]*(-5)+in_buf[371]*(-17)+in_buf[372]*(7)+in_buf[373]*(13)+in_buf[374]*(11)+in_buf[375]*(12)+in_buf[376]*(8)+in_buf[377]*(17)+in_buf[378]*(12)+in_buf[379]*(9)+in_buf[380]*(12)+in_buf[381]*(12)+in_buf[382]*(14)+in_buf[383]*(4)+in_buf[384]*(0)+in_buf[385]*(-3)+in_buf[386]*(-12)+in_buf[387]*(-6)+in_buf[388]*(-41)+in_buf[389]*(-45)+in_buf[390]*(-53)+in_buf[391]*(-18)+in_buf[392]*(-14)+in_buf[393]*(7)+in_buf[394]*(-12)+in_buf[395]*(6)+in_buf[396]*(14)+in_buf[397]*(22)+in_buf[398]*(-26)+in_buf[399]*(-20)+in_buf[400]*(6)+in_buf[401]*(11)+in_buf[402]*(-10)+in_buf[403]*(3)+in_buf[404]*(12)+in_buf[405]*(8)+in_buf[406]*(7)+in_buf[407]*(0)+in_buf[408]*(0)+in_buf[409]*(4)+in_buf[410]*(6)+in_buf[411]*(11)+in_buf[412]*(7)+in_buf[413]*(19)+in_buf[414]*(5)+in_buf[415]*(1)+in_buf[416]*(-16)+in_buf[417]*(-11)+in_buf[418]*(-30)+in_buf[419]*(-16)+in_buf[420]*(-12)+in_buf[421]*(11)+in_buf[422]*(32)+in_buf[423]*(15)+in_buf[424]*(22)+in_buf[425]*(-12)+in_buf[426]*(-27)+in_buf[427]*(-2)+in_buf[428]*(20)+in_buf[429]*(8)+in_buf[430]*(-1)+in_buf[431]*(5)+in_buf[432]*(5)+in_buf[433]*(15)+in_buf[434]*(15)+in_buf[435]*(6)+in_buf[436]*(15)+in_buf[437]*(0)+in_buf[438]*(-11)+in_buf[439]*(4)+in_buf[440]*(8)+in_buf[441]*(19)+in_buf[442]*(16)+in_buf[443]*(-7)+in_buf[444]*(-30)+in_buf[445]*(-11)+in_buf[446]*(13)+in_buf[447]*(-21)+in_buf[448]*(5)+in_buf[449]*(22)+in_buf[450]*(23)+in_buf[451]*(9)+in_buf[452]*(16)+in_buf[453]*(-21)+in_buf[454]*(-13)+in_buf[455]*(13)+in_buf[456]*(22)+in_buf[457]*(22)+in_buf[458]*(7)+in_buf[459]*(8)+in_buf[460]*(16)+in_buf[461]*(11)+in_buf[462]*(13)+in_buf[463]*(1)+in_buf[464]*(5)+in_buf[465]*(-12)+in_buf[466]*(4)+in_buf[467]*(0)+in_buf[468]*(11)+in_buf[469]*(14)+in_buf[470]*(-1)+in_buf[471]*(-2)+in_buf[472]*(-13)+in_buf[473]*(-25)+in_buf[474]*(-17)+in_buf[475]*(-27)+in_buf[476]*(0)+in_buf[477]*(10)+in_buf[478]*(23)+in_buf[479]*(13)+in_buf[480]*(31)+in_buf[481]*(-19)+in_buf[482]*(-31)+in_buf[483]*(3)+in_buf[484]*(12)+in_buf[485]*(2)+in_buf[486]*(-3)+in_buf[487]*(-8)+in_buf[488]*(8)+in_buf[489]*(14)+in_buf[490]*(3)+in_buf[491]*(-8)+in_buf[492]*(0)+in_buf[493]*(-9)+in_buf[494]*(1)+in_buf[495]*(7)+in_buf[496]*(-3)+in_buf[497]*(16)+in_buf[498]*(4)+in_buf[499]*(8)+in_buf[500]*(-23)+in_buf[501]*(-37)+in_buf[502]*(-12)+in_buf[503]*(-32)+in_buf[504]*(-28)+in_buf[505]*(11)+in_buf[506]*(24)+in_buf[507]*(16)+in_buf[508]*(21)+in_buf[509]*(-16)+in_buf[510]*(-16)+in_buf[511]*(-10)+in_buf[512]*(-9)+in_buf[513]*(2)+in_buf[514]*(-12)+in_buf[515]*(-1)+in_buf[516]*(8)+in_buf[517]*(4)+in_buf[518]*(-12)+in_buf[519]*(-10)+in_buf[520]*(0)+in_buf[521]*(1)+in_buf[522]*(0)+in_buf[523]*(3)+in_buf[524]*(6)+in_buf[525]*(15)+in_buf[526]*(5)+in_buf[527]*(-12)+in_buf[528]*(-42)+in_buf[529]*(-67)+in_buf[530]*(-2)+in_buf[531]*(9)+in_buf[532]*(22)+in_buf[533]*(-28)+in_buf[534]*(-7)+in_buf[535]*(21)+in_buf[536]*(8)+in_buf[537]*(3)+in_buf[538]*(-13)+in_buf[539]*(0)+in_buf[540]*(-7)+in_buf[541]*(-4)+in_buf[542]*(-3)+in_buf[543]*(-3)+in_buf[544]*(-17)+in_buf[545]*(-22)+in_buf[546]*(-8)+in_buf[547]*(-2)+in_buf[548]*(1)+in_buf[549]*(-2)+in_buf[550]*(3)+in_buf[551]*(9)+in_buf[552]*(5)+in_buf[553]*(11)+in_buf[554]*(-6)+in_buf[555]*(-27)+in_buf[556]*(-45)+in_buf[557]*(-52)+in_buf[558]*(-2)+in_buf[559]*(17)+in_buf[560]*(-1)+in_buf[561]*(0)+in_buf[562]*(-5)+in_buf[563]*(14)+in_buf[564]*(15)+in_buf[565]*(-10)+in_buf[566]*(-6)+in_buf[567]*(5)+in_buf[568]*(-9)+in_buf[569]*(-8)+in_buf[570]*(-3)+in_buf[571]*(-18)+in_buf[572]*(-20)+in_buf[573]*(-27)+in_buf[574]*(3)+in_buf[575]*(0)+in_buf[576]*(0)+in_buf[577]*(-6)+in_buf[578]*(9)+in_buf[579]*(5)+in_buf[580]*(13)+in_buf[581]*(2)+in_buf[582]*(-17)+in_buf[583]*(-29)+in_buf[584]*(-19)+in_buf[585]*(-31)+in_buf[586]*(-6)+in_buf[587]*(18)+in_buf[588]*(11)+in_buf[589]*(7)+in_buf[590]*(27)+in_buf[591]*(23)+in_buf[592]*(-9)+in_buf[593]*(-8)+in_buf[594]*(-1)+in_buf[595]*(-8)+in_buf[596]*(-2)+in_buf[597]*(-10)+in_buf[598]*(-2)+in_buf[599]*(-8)+in_buf[600]*(-11)+in_buf[601]*(-15)+in_buf[602]*(2)+in_buf[603]*(1)+in_buf[604]*(2)+in_buf[605]*(1)+in_buf[606]*(6)+in_buf[607]*(2)+in_buf[608]*(3)+in_buf[609]*(-3)+in_buf[610]*(-3)+in_buf[611]*(-12)+in_buf[612]*(-24)+in_buf[613]*(1)+in_buf[614]*(-31)+in_buf[615]*(-1)+in_buf[616]*(16)+in_buf[617]*(19)+in_buf[618]*(27)+in_buf[619]*(14)+in_buf[620]*(-6)+in_buf[621]*(-12)+in_buf[622]*(-10)+in_buf[623]*(-17)+in_buf[624]*(-13)+in_buf[625]*(-13)+in_buf[626]*(-6)+in_buf[627]*(0)+in_buf[628]*(-19)+in_buf[629]*(0)+in_buf[630]*(2)+in_buf[631]*(20)+in_buf[632]*(11)+in_buf[633]*(11)+in_buf[634]*(21)+in_buf[635]*(17)+in_buf[636]*(15)+in_buf[637]*(22)+in_buf[638]*(33)+in_buf[639]*(7)+in_buf[640]*(-26)+in_buf[641]*(10)+in_buf[642]*(14)+in_buf[643]*(-2)+in_buf[644]*(-3)+in_buf[645]*(0)+in_buf[646]*(25)+in_buf[647]*(0)+in_buf[648]*(-9)+in_buf[649]*(-8)+in_buf[650]*(-14)+in_buf[651]*(-8)+in_buf[652]*(-18)+in_buf[653]*(-4)+in_buf[654]*(3)+in_buf[655]*(0)+in_buf[656]*(4)+in_buf[657]*(11)+in_buf[658]*(9)+in_buf[659]*(19)+in_buf[660]*(13)+in_buf[661]*(25)+in_buf[662]*(32)+in_buf[663]*(15)+in_buf[664]*(12)+in_buf[665]*(17)+in_buf[666]*(6)+in_buf[667]*(0)+in_buf[668]*(-31)+in_buf[669]*(1)+in_buf[670]*(38)+in_buf[671]*(0)+in_buf[672]*(4)+in_buf[673]*(4)+in_buf[674]*(11)+in_buf[675]*(1)+in_buf[676]*(-11)+in_buf[677]*(-9)+in_buf[678]*(-6)+in_buf[679]*(0)+in_buf[680]*(0)+in_buf[681]*(-1)+in_buf[682]*(11)+in_buf[683]*(12)+in_buf[684]*(-4)+in_buf[685]*(-4)+in_buf[686]*(3)+in_buf[687]*(4)+in_buf[688]*(4)+in_buf[689]*(3)+in_buf[690]*(2)+in_buf[691]*(13)+in_buf[692]*(10)+in_buf[693]*(6)+in_buf[694]*(10)+in_buf[695]*(7)+in_buf[696]*(-22)+in_buf[697]*(4)+in_buf[698]*(-7)+in_buf[699]*(-3)+in_buf[700]*(2)+in_buf[701]*(3)+in_buf[702]*(28)+in_buf[703]*(-9)+in_buf[704]*(-31)+in_buf[705]*(-26)+in_buf[706]*(-27)+in_buf[707]*(-19)+in_buf[708]*(13)+in_buf[709]*(8)+in_buf[710]*(0)+in_buf[711]*(-10)+in_buf[712]*(1)+in_buf[713]*(-4)+in_buf[714]*(3)+in_buf[715]*(-16)+in_buf[716]*(-34)+in_buf[717]*(-14)+in_buf[718]*(6)+in_buf[719]*(-3)+in_buf[720]*(-4)+in_buf[721]*(-7)+in_buf[722]*(-16)+in_buf[723]*(-16)+in_buf[724]*(-24)+in_buf[725]*(-3)+in_buf[726]*(-13)+in_buf[727]*(2)+in_buf[728]*(4)+in_buf[729]*(-2)+in_buf[730]*(-2)+in_buf[731]*(-15)+in_buf[732]*(-24)+in_buf[733]*(-12)+in_buf[734]*(-17)+in_buf[735]*(-40)+in_buf[736]*(-43)+in_buf[737]*(-46)+in_buf[738]*(1)+in_buf[739]*(14)+in_buf[740]*(3)+in_buf[741]*(0)+in_buf[742]*(-1)+in_buf[743]*(-6)+in_buf[744]*(0)+in_buf[745]*(13)+in_buf[746]*(-7)+in_buf[747]*(-50)+in_buf[748]*(-32)+in_buf[749]*(-9)+in_buf[750]*(-20)+in_buf[751]*(-16)+in_buf[752]*(10)+in_buf[753]*(-4)+in_buf[754]*(-4)+in_buf[755]*(-1)+in_buf[756]*(4)+in_buf[757]*(-3)+in_buf[758]*(-2)+in_buf[759]*(0)+in_buf[760]*(-5)+in_buf[761]*(-9)+in_buf[762]*(-11)+in_buf[763]*(-10)+in_buf[764]*(-19)+in_buf[765]*(-28)+in_buf[766]*(-46)+in_buf[767]*(-34)+in_buf[768]*(-24)+in_buf[769]*(-46)+in_buf[770]*(-37)+in_buf[771]*(-3)+in_buf[772]*(-19)+in_buf[773]*(-25)+in_buf[774]*(2)+in_buf[775]*(14)+in_buf[776]*(20)+in_buf[777]*(3)+in_buf[778]*(6)+in_buf[779]*(16)+in_buf[780]*(-2)+in_buf[781]*(-1)+in_buf[782]*(-1)+in_buf[783]*(0);
assign in_buf_weight052=in_buf[0]*(-3)+in_buf[1]*(-3)+in_buf[2]*(0)+in_buf[3]*(-1)+in_buf[4]*(2)+in_buf[5]*(4)+in_buf[6]*(-2)+in_buf[7]*(-2)+in_buf[8]*(0)+in_buf[9]*(-2)+in_buf[10]*(3)+in_buf[11]*(-1)+in_buf[12]*(13)+in_buf[13]*(15)+in_buf[14]*(-2)+in_buf[15]*(0)+in_buf[16]*(-2)+in_buf[17]*(4)+in_buf[18]*(-1)+in_buf[19]*(0)+in_buf[20]*(3)+in_buf[21]*(4)+in_buf[22]*(-1)+in_buf[23]*(-2)+in_buf[24]*(-1)+in_buf[25]*(0)+in_buf[26]*(0)+in_buf[27]*(0)+in_buf[28]*(1)+in_buf[29]*(4)+in_buf[30]*(-2)+in_buf[31]*(2)+in_buf[32]*(6)+in_buf[33]*(4)+in_buf[34]*(11)+in_buf[35]*(8)+in_buf[36]*(9)+in_buf[37]*(15)+in_buf[38]*(17)+in_buf[39]*(9)+in_buf[40]*(28)+in_buf[41]*(46)+in_buf[42]*(54)+in_buf[43]*(56)+in_buf[44]*(35)+in_buf[45]*(39)+in_buf[46]*(24)+in_buf[47]*(17)+in_buf[48]*(13)+in_buf[49]*(0)+in_buf[50]*(6)+in_buf[51]*(7)+in_buf[52]*(-2)+in_buf[53]*(0)+in_buf[54]*(1)+in_buf[55]*(1)+in_buf[56]*(4)+in_buf[57]*(0)+in_buf[58]*(19)+in_buf[59]*(-5)+in_buf[60]*(8)+in_buf[61]*(8)+in_buf[62]*(18)+in_buf[63]*(13)+in_buf[64]*(-7)+in_buf[65]*(-25)+in_buf[66]*(-2)+in_buf[67]*(26)+in_buf[68]*(9)+in_buf[69]*(16)+in_buf[70]*(21)+in_buf[71]*(51)+in_buf[72]*(71)+in_buf[73]*(70)+in_buf[74]*(69)+in_buf[75]*(52)+in_buf[76]*(37)+in_buf[77]*(27)+in_buf[78]*(23)+in_buf[79]*(34)+in_buf[80]*(0)+in_buf[81]*(3)+in_buf[82]*(3)+in_buf[83]*(0)+in_buf[84]*(1)+in_buf[85]*(0)+in_buf[86]*(17)+in_buf[87]*(5)+in_buf[88]*(12)+in_buf[89]*(-16)+in_buf[90]*(14)+in_buf[91]*(19)+in_buf[92]*(0)+in_buf[93]*(5)+in_buf[94]*(21)+in_buf[95]*(-18)+in_buf[96]*(0)+in_buf[97]*(29)+in_buf[98]*(26)+in_buf[99]*(34)+in_buf[100]*(22)+in_buf[101]*(28)+in_buf[102]*(46)+in_buf[103]*(53)+in_buf[104]*(47)+in_buf[105]*(23)+in_buf[106]*(9)+in_buf[107]*(4)+in_buf[108]*(29)+in_buf[109]*(13)+in_buf[110]*(5)+in_buf[111]*(1)+in_buf[112]*(2)+in_buf[113]*(0)+in_buf[114]*(4)+in_buf[115]*(-12)+in_buf[116]*(-8)+in_buf[117]*(-4)+in_buf[118]*(12)+in_buf[119]*(-11)+in_buf[120]*(-20)+in_buf[121]*(-7)+in_buf[122]*(2)+in_buf[123]*(-9)+in_buf[124]*(-14)+in_buf[125]*(-14)+in_buf[126]*(-7)+in_buf[127]*(21)+in_buf[128]*(23)+in_buf[129]*(3)+in_buf[130]*(15)+in_buf[131]*(8)+in_buf[132]*(7)+in_buf[133]*(44)+in_buf[134]*(44)+in_buf[135]*(38)+in_buf[136]*(13)+in_buf[137]*(36)+in_buf[138]*(37)+in_buf[139]*(0)+in_buf[140]*(0)+in_buf[141]*(-3)+in_buf[142]*(9)+in_buf[143]*(-22)+in_buf[144]*(-16)+in_buf[145]*(16)+in_buf[146]*(1)+in_buf[147]*(-8)+in_buf[148]*(4)+in_buf[149]*(10)+in_buf[150]*(22)+in_buf[151]*(0)+in_buf[152]*(-4)+in_buf[153]*(-1)+in_buf[154]*(6)+in_buf[155]*(5)+in_buf[156]*(25)+in_buf[157]*(22)+in_buf[158]*(22)+in_buf[159]*(9)+in_buf[160]*(12)+in_buf[161]*(26)+in_buf[162]*(48)+in_buf[163]*(39)+in_buf[164]*(4)+in_buf[165]*(20)+in_buf[166]*(12)+in_buf[167]*(4)+in_buf[168]*(3)+in_buf[169]*(11)+in_buf[170]*(0)+in_buf[171]*(-56)+in_buf[172]*(-13)+in_buf[173]*(12)+in_buf[174]*(-5)+in_buf[175]*(19)+in_buf[176]*(21)+in_buf[177]*(17)+in_buf[178]*(11)+in_buf[179]*(23)+in_buf[180]*(17)+in_buf[181]*(9)+in_buf[182]*(14)+in_buf[183]*(17)+in_buf[184]*(17)+in_buf[185]*(24)+in_buf[186]*(39)+in_buf[187]*(30)+in_buf[188]*(27)+in_buf[189]*(27)+in_buf[190]*(29)+in_buf[191]*(-1)+in_buf[192]*(3)+in_buf[193]*(15)+in_buf[194]*(22)+in_buf[195]*(7)+in_buf[196]*(-4)+in_buf[197]*(20)+in_buf[198]*(-13)+in_buf[199]*(-57)+in_buf[200]*(-20)+in_buf[201]*(14)+in_buf[202]*(1)+in_buf[203]*(17)+in_buf[204]*(18)+in_buf[205]*(18)+in_buf[206]*(20)+in_buf[207]*(20)+in_buf[208]*(15)+in_buf[209]*(3)+in_buf[210]*(20)+in_buf[211]*(23)+in_buf[212]*(27)+in_buf[213]*(23)+in_buf[214]*(30)+in_buf[215]*(33)+in_buf[216]*(24)+in_buf[217]*(0)+in_buf[218]*(0)+in_buf[219]*(-8)+in_buf[220]*(-24)+in_buf[221]*(-3)+in_buf[222]*(22)+in_buf[223]*(7)+in_buf[224]*(-1)+in_buf[225]*(19)+in_buf[226]*(-28)+in_buf[227]*(-40)+in_buf[228]*(-29)+in_buf[229]*(-4)+in_buf[230]*(9)+in_buf[231]*(17)+in_buf[232]*(0)+in_buf[233]*(12)+in_buf[234]*(14)+in_buf[235]*(17)+in_buf[236]*(11)+in_buf[237]*(-5)+in_buf[238]*(-6)+in_buf[239]*(-13)+in_buf[240]*(-26)+in_buf[241]*(-27)+in_buf[242]*(-16)+in_buf[243]*(-16)+in_buf[244]*(-25)+in_buf[245]*(-25)+in_buf[246]*(-8)+in_buf[247]*(-15)+in_buf[248]*(-45)+in_buf[249]*(-29)+in_buf[250]*(17)+in_buf[251]*(4)+in_buf[252]*(3)+in_buf[253]*(19)+in_buf[254]*(-50)+in_buf[255]*(-51)+in_buf[256]*(-10)+in_buf[257]*(-6)+in_buf[258]*(8)+in_buf[259]*(7)+in_buf[260]*(16)+in_buf[261]*(6)+in_buf[262]*(0)+in_buf[263]*(9)+in_buf[264]*(0)+in_buf[265]*(-14)+in_buf[266]*(-32)+in_buf[267]*(-50)+in_buf[268]*(-79)+in_buf[269]*(-98)+in_buf[270]*(-83)+in_buf[271]*(-84)+in_buf[272]*(-70)+in_buf[273]*(-64)+in_buf[274]*(-40)+in_buf[275]*(-47)+in_buf[276]*(-41)+in_buf[277]*(-26)+in_buf[278]*(5)+in_buf[279]*(5)+in_buf[280]*(0)+in_buf[281]*(12)+in_buf[282]*(-27)+in_buf[283]*(-32)+in_buf[284]*(-10)+in_buf[285]*(0)+in_buf[286]*(-10)+in_buf[287]*(-2)+in_buf[288]*(12)+in_buf[289]*(-3)+in_buf[290]*(-11)+in_buf[291]*(0)+in_buf[292]*(-3)+in_buf[293]*(-15)+in_buf[294]*(-41)+in_buf[295]*(-44)+in_buf[296]*(-41)+in_buf[297]*(-63)+in_buf[298]*(-87)+in_buf[299]*(-90)+in_buf[300]*(-80)+in_buf[301]*(-90)+in_buf[302]*(-87)+in_buf[303]*(-100)+in_buf[304]*(-73)+in_buf[305]*(-29)+in_buf[306]*(1)+in_buf[307]*(11)+in_buf[308]*(-2)+in_buf[309]*(-16)+in_buf[310]*(-18)+in_buf[311]*(-29)+in_buf[312]*(-13)+in_buf[313]*(7)+in_buf[314]*(-7)+in_buf[315]*(-11)+in_buf[316]*(-6)+in_buf[317]*(-17)+in_buf[318]*(-9)+in_buf[319]*(-12)+in_buf[320]*(-11)+in_buf[321]*(-15)+in_buf[322]*(-19)+in_buf[323]*(-7)+in_buf[324]*(19)+in_buf[325]*(21)+in_buf[326]*(3)+in_buf[327]*(-25)+in_buf[328]*(-43)+in_buf[329]*(-53)+in_buf[330]*(-70)+in_buf[331]*(-98)+in_buf[332]*(-79)+in_buf[333]*(-47)+in_buf[334]*(-2)+in_buf[335]*(12)+in_buf[336]*(-3)+in_buf[337]*(-18)+in_buf[338]*(-25)+in_buf[339]*(-7)+in_buf[340]*(-13)+in_buf[341]*(10)+in_buf[342]*(6)+in_buf[343]*(-5)+in_buf[344]*(6)+in_buf[345]*(-19)+in_buf[346]*(4)+in_buf[347]*(-4)+in_buf[348]*(-11)+in_buf[349]*(-12)+in_buf[350]*(-8)+in_buf[351]*(6)+in_buf[352]*(18)+in_buf[353]*(10)+in_buf[354]*(30)+in_buf[355]*(0)+in_buf[356]*(-1)+in_buf[357]*(-9)+in_buf[358]*(-23)+in_buf[359]*(-40)+in_buf[360]*(-66)+in_buf[361]*(-40)+in_buf[362]*(0)+in_buf[363]*(17)+in_buf[364]*(-3)+in_buf[365]*(-5)+in_buf[366]*(-9)+in_buf[367]*(-9)+in_buf[368]*(14)+in_buf[369]*(14)+in_buf[370]*(20)+in_buf[371]*(15)+in_buf[372]*(-9)+in_buf[373]*(-7)+in_buf[374]*(0)+in_buf[375]*(-11)+in_buf[376]*(-4)+in_buf[377]*(-9)+in_buf[378]*(-3)+in_buf[379]*(8)+in_buf[380]*(-7)+in_buf[381]*(6)+in_buf[382]*(6)+in_buf[383]*(12)+in_buf[384]*(17)+in_buf[385]*(-1)+in_buf[386]*(-10)+in_buf[387]*(-7)+in_buf[388]*(0)+in_buf[389]*(-42)+in_buf[390]*(-3)+in_buf[391]*(-16)+in_buf[392]*(15)+in_buf[393]*(1)+in_buf[394]*(-6)+in_buf[395]*(1)+in_buf[396]*(13)+in_buf[397]*(0)+in_buf[398]*(22)+in_buf[399]*(13)+in_buf[400]*(14)+in_buf[401]*(-7)+in_buf[402]*(7)+in_buf[403]*(-7)+in_buf[404]*(-21)+in_buf[405]*(-18)+in_buf[406]*(7)+in_buf[407]*(9)+in_buf[408]*(3)+in_buf[409]*(1)+in_buf[410]*(14)+in_buf[411]*(10)+in_buf[412]*(16)+in_buf[413]*(3)+in_buf[414]*(2)+in_buf[415]*(9)+in_buf[416]*(36)+in_buf[417]*(-15)+in_buf[418]*(-21)+in_buf[419]*(-17)+in_buf[420]*(16)+in_buf[421]*(9)+in_buf[422]*(17)+in_buf[423]*(-6)+in_buf[424]*(-42)+in_buf[425]*(-17)+in_buf[426]*(-9)+in_buf[427]*(-3)+in_buf[428]*(0)+in_buf[429]*(5)+in_buf[430]*(2)+in_buf[431]*(-7)+in_buf[432]*(-15)+in_buf[433]*(-19)+in_buf[434]*(6)+in_buf[435]*(11)+in_buf[436]*(4)+in_buf[437]*(8)+in_buf[438]*(19)+in_buf[439]*(4)+in_buf[440]*(15)+in_buf[441]*(25)+in_buf[442]*(4)+in_buf[443]*(16)+in_buf[444]*(37)+in_buf[445]*(14)+in_buf[446]*(-4)+in_buf[447]*(-16)+in_buf[448]*(0)+in_buf[449]*(4)+in_buf[450]*(15)+in_buf[451]*(9)+in_buf[452]*(-54)+in_buf[453]*(-43)+in_buf[454]*(-47)+in_buf[455]*(-23)+in_buf[456]*(-22)+in_buf[457]*(-11)+in_buf[458]*(-6)+in_buf[459]*(-1)+in_buf[460]*(-26)+in_buf[461]*(-10)+in_buf[462]*(11)+in_buf[463]*(16)+in_buf[464]*(0)+in_buf[465]*(-1)+in_buf[466]*(6)+in_buf[467]*(11)+in_buf[468]*(22)+in_buf[469]*(16)+in_buf[470]*(21)+in_buf[471]*(8)+in_buf[472]*(36)+in_buf[473]*(34)+in_buf[474]*(8)+in_buf[475]*(-21)+in_buf[476]*(-3)+in_buf[477]*(-1)+in_buf[478]*(-19)+in_buf[479]*(22)+in_buf[480]*(-40)+in_buf[481]*(-45)+in_buf[482]*(-36)+in_buf[483]*(-21)+in_buf[484]*(-13)+in_buf[485]*(-18)+in_buf[486]*(-14)+in_buf[487]*(-6)+in_buf[488]*(-25)+in_buf[489]*(-25)+in_buf[490]*(9)+in_buf[491]*(9)+in_buf[492]*(-9)+in_buf[493]*(-8)+in_buf[494]*(5)+in_buf[495]*(7)+in_buf[496]*(5)+in_buf[497]*(20)+in_buf[498]*(11)+in_buf[499]*(6)+in_buf[500]*(17)+in_buf[501]*(-18)+in_buf[502]*(-31)+in_buf[503]*(-36)+in_buf[504]*(-2)+in_buf[505]*(-13)+in_buf[506]*(-27)+in_buf[507]*(28)+in_buf[508]*(4)+in_buf[509]*(-18)+in_buf[510]*(-17)+in_buf[511]*(-17)+in_buf[512]*(-6)+in_buf[513]*(-10)+in_buf[514]*(-16)+in_buf[515]*(-26)+in_buf[516]*(-38)+in_buf[517]*(-31)+in_buf[518]*(11)+in_buf[519]*(16)+in_buf[520]*(12)+in_buf[521]*(11)+in_buf[522]*(5)+in_buf[523]*(-6)+in_buf[524]*(15)+in_buf[525]*(24)+in_buf[526]*(4)+in_buf[527]*(0)+in_buf[528]*(15)+in_buf[529]*(-33)+in_buf[530]*(-38)+in_buf[531]*(-41)+in_buf[532]*(-1)+in_buf[533]*(-38)+in_buf[534]*(13)+in_buf[535]*(26)+in_buf[536]*(17)+in_buf[537]*(-7)+in_buf[538]*(-9)+in_buf[539]*(-23)+in_buf[540]*(-16)+in_buf[541]*(-8)+in_buf[542]*(-11)+in_buf[543]*(6)+in_buf[544]*(-6)+in_buf[545]*(-18)+in_buf[546]*(7)+in_buf[547]*(19)+in_buf[548]*(23)+in_buf[549]*(9)+in_buf[550]*(10)+in_buf[551]*(4)+in_buf[552]*(21)+in_buf[553]*(22)+in_buf[554]*(13)+in_buf[555]*(9)+in_buf[556]*(26)+in_buf[557]*(5)+in_buf[558]*(-41)+in_buf[559]*(-27)+in_buf[560]*(0)+in_buf[561]*(-19)+in_buf[562]*(11)+in_buf[563]*(34)+in_buf[564]*(41)+in_buf[565]*(3)+in_buf[566]*(-13)+in_buf[567]*(-19)+in_buf[568]*(-11)+in_buf[569]*(0)+in_buf[570]*(-3)+in_buf[571]*(12)+in_buf[572]*(-5)+in_buf[573]*(-8)+in_buf[574]*(9)+in_buf[575]*(22)+in_buf[576]*(25)+in_buf[577]*(27)+in_buf[578]*(16)+in_buf[579]*(9)+in_buf[580]*(2)+in_buf[581]*(8)+in_buf[582]*(28)+in_buf[583]*(19)+in_buf[584]*(11)+in_buf[585]*(32)+in_buf[586]*(-13)+in_buf[587]*(3)+in_buf[588]*(-1)+in_buf[589]*(-20)+in_buf[590]*(-39)+in_buf[591]*(19)+in_buf[592]*(42)+in_buf[593]*(22)+in_buf[594]*(4)+in_buf[595]*(12)+in_buf[596]*(3)+in_buf[597]*(1)+in_buf[598]*(14)+in_buf[599]*(18)+in_buf[600]*(20)+in_buf[601]*(9)+in_buf[602]*(18)+in_buf[603]*(28)+in_buf[604]*(16)+in_buf[605]*(12)+in_buf[606]*(14)+in_buf[607]*(3)+in_buf[608]*(11)+in_buf[609]*(25)+in_buf[610]*(11)+in_buf[611]*(-1)+in_buf[612]*(25)+in_buf[613]*(28)+in_buf[614]*(20)+in_buf[615]*(-3)+in_buf[616]*(-1)+in_buf[617]*(-29)+in_buf[618]*(-15)+in_buf[619]*(6)+in_buf[620]*(12)+in_buf[621]*(16)+in_buf[622]*(0)+in_buf[623]*(-1)+in_buf[624]*(11)+in_buf[625]*(4)+in_buf[626]*(0)+in_buf[627]*(8)+in_buf[628]*(7)+in_buf[629]*(2)+in_buf[630]*(8)+in_buf[631]*(16)+in_buf[632]*(13)+in_buf[633]*(9)+in_buf[634]*(-1)+in_buf[635]*(9)+in_buf[636]*(18)+in_buf[637]*(8)+in_buf[638]*(2)+in_buf[639]*(6)+in_buf[640]*(13)+in_buf[641]*(27)+in_buf[642]*(22)+in_buf[643]*(-5)+in_buf[644]*(3)+in_buf[645]*(-2)+in_buf[646]*(19)+in_buf[647]*(27)+in_buf[648]*(24)+in_buf[649]*(15)+in_buf[650]*(20)+in_buf[651]*(3)+in_buf[652]*(10)+in_buf[653]*(11)+in_buf[654]*(9)+in_buf[655]*(7)+in_buf[656]*(11)+in_buf[657]*(10)+in_buf[658]*(11)+in_buf[659]*(7)+in_buf[660]*(1)+in_buf[661]*(10)+in_buf[662]*(0)+in_buf[663]*(3)+in_buf[664]*(12)+in_buf[665]*(3)+in_buf[666]*(9)+in_buf[667]*(-5)+in_buf[668]*(12)+in_buf[669]*(17)+in_buf[670]*(30)+in_buf[671]*(0)+in_buf[672]*(1)+in_buf[673]*(2)+in_buf[674]*(-13)+in_buf[675]*(17)+in_buf[676]*(20)+in_buf[677]*(12)+in_buf[678]*(37)+in_buf[679]*(54)+in_buf[680]*(33)+in_buf[681]*(34)+in_buf[682]*(17)+in_buf[683]*(15)+in_buf[684]*(24)+in_buf[685]*(18)+in_buf[686]*(14)+in_buf[687]*(10)+in_buf[688]*(3)+in_buf[689]*(13)+in_buf[690]*(21)+in_buf[691]*(-9)+in_buf[692]*(9)+in_buf[693]*(9)+in_buf[694]*(-1)+in_buf[695]*(-34)+in_buf[696]*(-12)+in_buf[697]*(-4)+in_buf[698]*(2)+in_buf[699]*(0)+in_buf[700]*(-2)+in_buf[701]*(2)+in_buf[702]*(8)+in_buf[703]*(11)+in_buf[704]*(4)+in_buf[705]*(-1)+in_buf[706]*(27)+in_buf[707]*(42)+in_buf[708]*(27)+in_buf[709]*(39)+in_buf[710]*(23)+in_buf[711]*(34)+in_buf[712]*(42)+in_buf[713]*(30)+in_buf[714]*(1)+in_buf[715]*(9)+in_buf[716]*(2)+in_buf[717]*(-14)+in_buf[718]*(-13)+in_buf[719]*(38)+in_buf[720]*(32)+in_buf[721]*(22)+in_buf[722]*(24)+in_buf[723]*(-7)+in_buf[724]*(12)+in_buf[725]*(4)+in_buf[726]*(-1)+in_buf[727]*(-2)+in_buf[728]*(1)+in_buf[729]*(-3)+in_buf[730]*(-1)+in_buf[731]*(2)+in_buf[732]*(-4)+in_buf[733]*(-6)+in_buf[734]*(-5)+in_buf[735]*(-27)+in_buf[736]*(-41)+in_buf[737]*(-20)+in_buf[738]*(15)+in_buf[739]*(1)+in_buf[740]*(-24)+in_buf[741]*(12)+in_buf[742]*(0)+in_buf[743]*(-10)+in_buf[744]*(-45)+in_buf[745]*(-51)+in_buf[746]*(-1)+in_buf[747]*(21)+in_buf[748]*(33)+in_buf[749]*(34)+in_buf[750]*(36)+in_buf[751]*(2)+in_buf[752]*(-2)+in_buf[753]*(4)+in_buf[754]*(0)+in_buf[755]*(3)+in_buf[756]*(0)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(0)+in_buf[760]*(2)+in_buf[761]*(3)+in_buf[762]*(-1)+in_buf[763]*(2)+in_buf[764]*(-1)+in_buf[765]*(0)+in_buf[766]*(-11)+in_buf[767]*(-4)+in_buf[768]*(-6)+in_buf[769]*(-8)+in_buf[770]*(-10)+in_buf[771]*(-7)+in_buf[772]*(-1)+in_buf[773]*(2)+in_buf[774]*(-2)+in_buf[775]*(-15)+in_buf[776]*(-18)+in_buf[777]*(24)+in_buf[778]*(19)+in_buf[779]*(-2)+in_buf[780]*(4)+in_buf[781]*(0)+in_buf[782]*(0)+in_buf[783]*(-4);
assign in_buf_weight053=in_buf[0]*(3)+in_buf[1]*(2)+in_buf[2]*(-2)+in_buf[3]*(-2)+in_buf[4]*(3)+in_buf[5]*(0)+in_buf[6]*(-1)+in_buf[7]*(3)+in_buf[8]*(0)+in_buf[9]*(2)+in_buf[10]*(-3)+in_buf[11]*(0)+in_buf[12]*(17)+in_buf[13]*(12)+in_buf[14]*(1)+in_buf[15]*(-5)+in_buf[16]*(0)+in_buf[17]*(0)+in_buf[18]*(0)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(2)+in_buf[22]*(-1)+in_buf[23]*(3)+in_buf[24]*(-1)+in_buf[25]*(3)+in_buf[26]*(2)+in_buf[27]*(-2)+in_buf[28]*(-1)+in_buf[29]*(-1)+in_buf[30]*(2)+in_buf[31]*(2)+in_buf[32]*(2)+in_buf[33]*(5)+in_buf[34]*(7)+in_buf[35]*(10)+in_buf[36]*(14)+in_buf[37]*(11)+in_buf[38]*(24)+in_buf[39]*(4)+in_buf[40]*(2)+in_buf[41]*(12)+in_buf[42]*(25)+in_buf[43]*(18)+in_buf[44]*(-2)+in_buf[45]*(-2)+in_buf[46]*(21)+in_buf[47]*(19)+in_buf[48]*(17)+in_buf[49]*(12)+in_buf[50]*(6)+in_buf[51]*(10)+in_buf[52]*(2)+in_buf[53]*(-2)+in_buf[54]*(-2)+in_buf[55]*(-1)+in_buf[56]*(4)+in_buf[57]*(2)+in_buf[58]*(3)+in_buf[59]*(0)+in_buf[60]*(1)+in_buf[61]*(8)+in_buf[62]*(21)+in_buf[63]*(18)+in_buf[64]*(36)+in_buf[65]*(27)+in_buf[66]*(16)+in_buf[67]*(45)+in_buf[68]*(36)+in_buf[69]*(34)+in_buf[70]*(58)+in_buf[71]*(52)+in_buf[72]*(6)+in_buf[73]*(1)+in_buf[74]*(14)+in_buf[75]*(7)+in_buf[76]*(14)+in_buf[77]*(6)+in_buf[78]*(9)+in_buf[79]*(16)+in_buf[80]*(17)+in_buf[81]*(3)+in_buf[82]*(1)+in_buf[83]*(4)+in_buf[84]*(2)+in_buf[85]*(0)+in_buf[86]*(-17)+in_buf[87]*(0)+in_buf[88]*(12)+in_buf[89]*(17)+in_buf[90]*(46)+in_buf[91]*(27)+in_buf[92]*(10)+in_buf[93]*(24)+in_buf[94]*(20)+in_buf[95]*(-5)+in_buf[96]*(-13)+in_buf[97]*(-10)+in_buf[98]*(-20)+in_buf[99]*(-22)+in_buf[100]*(-15)+in_buf[101]*(-6)+in_buf[102]*(-15)+in_buf[103]*(29)+in_buf[104]*(3)+in_buf[105]*(-8)+in_buf[106]*(-1)+in_buf[107]*(6)+in_buf[108]*(21)+in_buf[109]*(-2)+in_buf[110]*(2)+in_buf[111]*(1)+in_buf[112]*(0)+in_buf[113]*(4)+in_buf[114]*(-5)+in_buf[115]*(-9)+in_buf[116]*(34)+in_buf[117]*(50)+in_buf[118]*(31)+in_buf[119]*(20)+in_buf[120]*(29)+in_buf[121]*(16)+in_buf[122]*(15)+in_buf[123]*(-11)+in_buf[124]*(-18)+in_buf[125]*(-22)+in_buf[126]*(-26)+in_buf[127]*(-36)+in_buf[128]*(0)+in_buf[129]*(3)+in_buf[130]*(5)+in_buf[131]*(26)+in_buf[132]*(-4)+in_buf[133]*(-10)+in_buf[134]*(-6)+in_buf[135]*(-5)+in_buf[136]*(3)+in_buf[137]*(6)+in_buf[138]*(19)+in_buf[139]*(2)+in_buf[140]*(-2)+in_buf[141]*(2)+in_buf[142]*(6)+in_buf[143]*(21)+in_buf[144]*(47)+in_buf[145]*(53)+in_buf[146]*(31)+in_buf[147]*(28)+in_buf[148]*(35)+in_buf[149]*(6)+in_buf[150]*(-5)+in_buf[151]*(-11)+in_buf[152]*(7)+in_buf[153]*(-11)+in_buf[154]*(-18)+in_buf[155]*(-27)+in_buf[156]*(-6)+in_buf[157]*(-16)+in_buf[158]*(-11)+in_buf[159]*(-10)+in_buf[160]*(-23)+in_buf[161]*(-17)+in_buf[162]*(-17)+in_buf[163]*(-8)+in_buf[164]*(0)+in_buf[165]*(15)+in_buf[166]*(19)+in_buf[167]*(8)+in_buf[168]*(-2)+in_buf[169]*(2)+in_buf[170]*(-2)+in_buf[171]*(27)+in_buf[172]*(23)+in_buf[173]*(18)+in_buf[174]*(17)+in_buf[175]*(10)+in_buf[176]*(10)+in_buf[177]*(10)+in_buf[178]*(-5)+in_buf[179]*(9)+in_buf[180]*(18)+in_buf[181]*(-4)+in_buf[182]*(-11)+in_buf[183]*(-20)+in_buf[184]*(-17)+in_buf[185]*(0)+in_buf[186]*(0)+in_buf[187]*(6)+in_buf[188]*(9)+in_buf[189]*(13)+in_buf[190]*(-19)+in_buf[191]*(8)+in_buf[192]*(-16)+in_buf[193]*(-11)+in_buf[194]*(-11)+in_buf[195]*(-19)+in_buf[196]*(0)+in_buf[197]*(9)+in_buf[198]*(26)+in_buf[199]*(31)+in_buf[200]*(20)+in_buf[201]*(-6)+in_buf[202]*(-2)+in_buf[203]*(8)+in_buf[204]*(0)+in_buf[205]*(9)+in_buf[206]*(1)+in_buf[207]*(9)+in_buf[208]*(7)+in_buf[209]*(-3)+in_buf[210]*(-12)+in_buf[211]*(-14)+in_buf[212]*(-18)+in_buf[213]*(1)+in_buf[214]*(20)+in_buf[215]*(6)+in_buf[216]*(8)+in_buf[217]*(20)+in_buf[218]*(9)+in_buf[219]*(11)+in_buf[220]*(-38)+in_buf[221]*(-26)+in_buf[222]*(-31)+in_buf[223]*(-23)+in_buf[224]*(-5)+in_buf[225]*(20)+in_buf[226]*(28)+in_buf[227]*(29)+in_buf[228]*(33)+in_buf[229]*(12)+in_buf[230]*(2)+in_buf[231]*(17)+in_buf[232]*(6)+in_buf[233]*(10)+in_buf[234]*(9)+in_buf[235]*(2)+in_buf[236]*(5)+in_buf[237]*(0)+in_buf[238]*(-2)+in_buf[239]*(-9)+in_buf[240]*(-17)+in_buf[241]*(-12)+in_buf[242]*(11)+in_buf[243]*(0)+in_buf[244]*(18)+in_buf[245]*(10)+in_buf[246]*(9)+in_buf[247]*(17)+in_buf[248]*(-45)+in_buf[249]*(-37)+in_buf[250]*(-3)+in_buf[251]*(-14)+in_buf[252]*(8)+in_buf[253]*(22)+in_buf[254]*(17)+in_buf[255]*(29)+in_buf[256]*(25)+in_buf[257]*(27)+in_buf[258]*(-3)+in_buf[259]*(6)+in_buf[260]*(8)+in_buf[261]*(5)+in_buf[262]*(-6)+in_buf[263]*(0)+in_buf[264]*(0)+in_buf[265]*(0)+in_buf[266]*(9)+in_buf[267]*(-7)+in_buf[268]*(-5)+in_buf[269]*(1)+in_buf[270]*(-1)+in_buf[271]*(-5)+in_buf[272]*(20)+in_buf[273]*(9)+in_buf[274]*(6)+in_buf[275]*(10)+in_buf[276]*(-27)+in_buf[277]*(-27)+in_buf[278]*(-15)+in_buf[279]*(-1)+in_buf[280]*(17)+in_buf[281]*(16)+in_buf[282]*(27)+in_buf[283]*(-6)+in_buf[284]*(23)+in_buf[285]*(19)+in_buf[286]*(12)+in_buf[287]*(11)+in_buf[288]*(7)+in_buf[289]*(3)+in_buf[290]*(8)+in_buf[291]*(7)+in_buf[292]*(-6)+in_buf[293]*(-3)+in_buf[294]*(-11)+in_buf[295]*(-7)+in_buf[296]*(4)+in_buf[297]*(3)+in_buf[298]*(-11)+in_buf[299]*(-8)+in_buf[300]*(-3)+in_buf[301]*(-5)+in_buf[302]*(-1)+in_buf[303]*(0)+in_buf[304]*(-2)+in_buf[305]*(-35)+in_buf[306]*(-43)+in_buf[307]*(-3)+in_buf[308]*(12)+in_buf[309]*(34)+in_buf[310]*(21)+in_buf[311]*(19)+in_buf[312]*(31)+in_buf[313]*(12)+in_buf[314]*(7)+in_buf[315]*(7)+in_buf[316]*(1)+in_buf[317]*(8)+in_buf[318]*(10)+in_buf[319]*(2)+in_buf[320]*(-8)+in_buf[321]*(-33)+in_buf[322]*(-24)+in_buf[323]*(-5)+in_buf[324]*(2)+in_buf[325]*(-10)+in_buf[326]*(0)+in_buf[327]*(-4)+in_buf[328]*(-8)+in_buf[329]*(-14)+in_buf[330]*(-7)+in_buf[331]*(-12)+in_buf[332]*(-18)+in_buf[333]*(-28)+in_buf[334]*(-26)+in_buf[335]*(-11)+in_buf[336]*(14)+in_buf[337]*(24)+in_buf[338]*(1)+in_buf[339]*(31)+in_buf[340]*(28)+in_buf[341]*(13)+in_buf[342]*(-21)+in_buf[343]*(2)+in_buf[344]*(1)+in_buf[345]*(-8)+in_buf[346]*(0)+in_buf[347]*(-2)+in_buf[348]*(-15)+in_buf[349]*(-26)+in_buf[350]*(-13)+in_buf[351]*(7)+in_buf[352]*(3)+in_buf[353]*(-4)+in_buf[354]*(1)+in_buf[355]*(-3)+in_buf[356]*(-1)+in_buf[357]*(-8)+in_buf[358]*(-10)+in_buf[359]*(-24)+in_buf[360]*(18)+in_buf[361]*(-6)+in_buf[362]*(-21)+in_buf[363]*(-2)+in_buf[364]*(-1)+in_buf[365]*(13)+in_buf[366]*(34)+in_buf[367]*(39)+in_buf[368]*(17)+in_buf[369]*(10)+in_buf[370]*(-3)+in_buf[371]*(1)+in_buf[372]*(-1)+in_buf[373]*(-2)+in_buf[374]*(-5)+in_buf[375]*(-10)+in_buf[376]*(-39)+in_buf[377]*(-28)+in_buf[378]*(-5)+in_buf[379]*(13)+in_buf[380]*(3)+in_buf[381]*(0)+in_buf[382]*(1)+in_buf[383]*(0)+in_buf[384]*(3)+in_buf[385]*(8)+in_buf[386]*(-2)+in_buf[387]*(-5)+in_buf[388]*(16)+in_buf[389]*(0)+in_buf[390]*(18)+in_buf[391]*(-7)+in_buf[392]*(-13)+in_buf[393]*(19)+in_buf[394]*(36)+in_buf[395]*(8)+in_buf[396]*(-3)+in_buf[397]*(23)+in_buf[398]*(8)+in_buf[399]*(-1)+in_buf[400]*(-4)+in_buf[401]*(-7)+in_buf[402]*(-2)+in_buf[403]*(-6)+in_buf[404]*(-16)+in_buf[405]*(-8)+in_buf[406]*(13)+in_buf[407]*(18)+in_buf[408]*(1)+in_buf[409]*(-1)+in_buf[410]*(2)+in_buf[411]*(28)+in_buf[412]*(5)+in_buf[413]*(8)+in_buf[414]*(21)+in_buf[415]*(22)+in_buf[416]*(5)+in_buf[417]*(-7)+in_buf[418]*(-1)+in_buf[419]*(0)+in_buf[420]*(-10)+in_buf[421]*(-9)+in_buf[422]*(28)+in_buf[423]*(1)+in_buf[424]*(-18)+in_buf[425]*(7)+in_buf[426]*(33)+in_buf[427]*(17)+in_buf[428]*(-13)+in_buf[429]*(-21)+in_buf[430]*(-24)+in_buf[431]*(-26)+in_buf[432]*(-29)+in_buf[433]*(21)+in_buf[434]*(44)+in_buf[435]*(21)+in_buf[436]*(4)+in_buf[437]*(11)+in_buf[438]*(2)+in_buf[439]*(21)+in_buf[440]*(15)+in_buf[441]*(0)+in_buf[442]*(18)+in_buf[443]*(12)+in_buf[444]*(-5)+in_buf[445]*(-3)+in_buf[446]*(-25)+in_buf[447]*(0)+in_buf[448]*(9)+in_buf[449]*(-5)+in_buf[450]*(24)+in_buf[451]*(2)+in_buf[452]*(-2)+in_buf[453]*(7)+in_buf[454]*(38)+in_buf[455]*(7)+in_buf[456]*(-16)+in_buf[457]*(-27)+in_buf[458]*(-43)+in_buf[459]*(-44)+in_buf[460]*(-17)+in_buf[461]*(23)+in_buf[462]*(48)+in_buf[463]*(24)+in_buf[464]*(21)+in_buf[465]*(18)+in_buf[466]*(15)+in_buf[467]*(22)+in_buf[468]*(3)+in_buf[469]*(17)+in_buf[470]*(14)+in_buf[471]*(-3)+in_buf[472]*(2)+in_buf[473]*(-23)+in_buf[474]*(-44)+in_buf[475]*(-5)+in_buf[476]*(2)+in_buf[477]*(5)+in_buf[478]*(23)+in_buf[479]*(-3)+in_buf[480]*(8)+in_buf[481]*(-2)+in_buf[482]*(-2)+in_buf[483]*(-40)+in_buf[484]*(-50)+in_buf[485]*(-67)+in_buf[486]*(-67)+in_buf[487]*(-22)+in_buf[488]*(18)+in_buf[489]*(45)+in_buf[490]*(46)+in_buf[491]*(19)+in_buf[492]*(17)+in_buf[493]*(24)+in_buf[494]*(21)+in_buf[495]*(5)+in_buf[496]*(13)+in_buf[497]*(10)+in_buf[498]*(23)+in_buf[499]*(9)+in_buf[500]*(21)+in_buf[501]*(0)+in_buf[502]*(-2)+in_buf[503]*(-3)+in_buf[504]*(21)+in_buf[505]*(10)+in_buf[506]*(25)+in_buf[507]*(20)+in_buf[508]*(1)+in_buf[509]*(-5)+in_buf[510]*(-28)+in_buf[511]*(-41)+in_buf[512]*(-57)+in_buf[513]*(-54)+in_buf[514]*(-57)+in_buf[515]*(-14)+in_buf[516]*(42)+in_buf[517]*(48)+in_buf[518]*(35)+in_buf[519]*(21)+in_buf[520]*(15)+in_buf[521]*(21)+in_buf[522]*(25)+in_buf[523]*(3)+in_buf[524]*(5)+in_buf[525]*(0)+in_buf[526]*(7)+in_buf[527]*(-23)+in_buf[528]*(-9)+in_buf[529]*(-16)+in_buf[530]*(25)+in_buf[531]*(7)+in_buf[532]*(-4)+in_buf[533]*(25)+in_buf[534]*(30)+in_buf[535]*(9)+in_buf[536]*(0)+in_buf[537]*(-29)+in_buf[538]*(-27)+in_buf[539]*(-51)+in_buf[540]*(-55)+in_buf[541]*(-42)+in_buf[542]*(-20)+in_buf[543]*(5)+in_buf[544]*(24)+in_buf[545]*(31)+in_buf[546]*(23)+in_buf[547]*(17)+in_buf[548]*(11)+in_buf[549]*(16)+in_buf[550]*(-4)+in_buf[551]*(-2)+in_buf[552]*(3)+in_buf[553]*(-16)+in_buf[554]*(-29)+in_buf[555]*(-43)+in_buf[556]*(-24)+in_buf[557]*(-43)+in_buf[558]*(20)+in_buf[559]*(4)+in_buf[560]*(0)+in_buf[561]*(0)+in_buf[562]*(15)+in_buf[563]*(-1)+in_buf[564]*(-41)+in_buf[565]*(-43)+in_buf[566]*(-24)+in_buf[567]*(-19)+in_buf[568]*(-31)+in_buf[569]*(-23)+in_buf[570]*(-4)+in_buf[571]*(6)+in_buf[572]*(22)+in_buf[573]*(14)+in_buf[574]*(19)+in_buf[575]*(21)+in_buf[576]*(14)+in_buf[577]*(9)+in_buf[578]*(-4)+in_buf[579]*(-8)+in_buf[580]*(-11)+in_buf[581]*(-37)+in_buf[582]*(-35)+in_buf[583]*(-47)+in_buf[584]*(-4)+in_buf[585]*(-29)+in_buf[586]*(17)+in_buf[587]*(6)+in_buf[588]*(-7)+in_buf[589]*(2)+in_buf[590]*(8)+in_buf[591]*(-12)+in_buf[592]*(-43)+in_buf[593]*(-44)+in_buf[594]*(-18)+in_buf[595]*(-41)+in_buf[596]*(-33)+in_buf[597]*(-21)+in_buf[598]*(0)+in_buf[599]*(-9)+in_buf[600]*(0)+in_buf[601]*(12)+in_buf[602]*(19)+in_buf[603]*(22)+in_buf[604]*(12)+in_buf[605]*(14)+in_buf[606]*(1)+in_buf[607]*(0)+in_buf[608]*(-24)+in_buf[609]*(-41)+in_buf[610]*(-25)+in_buf[611]*(-23)+in_buf[612]*(0)+in_buf[613]*(-2)+in_buf[614]*(0)+in_buf[615]*(0)+in_buf[616]*(-1)+in_buf[617]*(-4)+in_buf[618]*(3)+in_buf[619]*(-21)+in_buf[620]*(-23)+in_buf[621]*(-37)+in_buf[622]*(-40)+in_buf[623]*(-33)+in_buf[624]*(-28)+in_buf[625]*(-20)+in_buf[626]*(-20)+in_buf[627]*(-14)+in_buf[628]*(-16)+in_buf[629]*(3)+in_buf[630]*(2)+in_buf[631]*(6)+in_buf[632]*(12)+in_buf[633]*(10)+in_buf[634]*(0)+in_buf[635]*(-1)+in_buf[636]*(-32)+in_buf[637]*(-21)+in_buf[638]*(-5)+in_buf[639]*(0)+in_buf[640]*(0)+in_buf[641]*(14)+in_buf[642]*(19)+in_buf[643]*(2)+in_buf[644]*(0)+in_buf[645]*(2)+in_buf[646]*(-5)+in_buf[647]*(-37)+in_buf[648]*(-18)+in_buf[649]*(-22)+in_buf[650]*(-18)+in_buf[651]*(-20)+in_buf[652]*(-27)+in_buf[653]*(-12)+in_buf[654]*(-18)+in_buf[655]*(-15)+in_buf[656]*(-4)+in_buf[657]*(5)+in_buf[658]*(0)+in_buf[659]*(5)+in_buf[660]*(8)+in_buf[661]*(10)+in_buf[662]*(-2)+in_buf[663]*(-2)+in_buf[664]*(-18)+in_buf[665]*(0)+in_buf[666]*(11)+in_buf[667]*(7)+in_buf[668]*(1)+in_buf[669]*(10)+in_buf[670]*(12)+in_buf[671]*(-2)+in_buf[672]*(-3)+in_buf[673]*(3)+in_buf[674]*(9)+in_buf[675]*(-16)+in_buf[676]*(3)+in_buf[677]*(-3)+in_buf[678]*(-3)+in_buf[679]*(-16)+in_buf[680]*(-8)+in_buf[681]*(-6)+in_buf[682]*(-12)+in_buf[683]*(-7)+in_buf[684]*(-3)+in_buf[685]*(-5)+in_buf[686]*(9)+in_buf[687]*(5)+in_buf[688]*(2)+in_buf[689]*(0)+in_buf[690]*(1)+in_buf[691]*(6)+in_buf[692]*(9)+in_buf[693]*(-3)+in_buf[694]*(19)+in_buf[695]*(0)+in_buf[696]*(12)+in_buf[697]*(0)+in_buf[698]*(1)+in_buf[699]*(-3)+in_buf[700]*(0)+in_buf[701]*(2)+in_buf[702]*(-29)+in_buf[703]*(3)+in_buf[704]*(7)+in_buf[705]*(-27)+in_buf[706]*(6)+in_buf[707]*(0)+in_buf[708]*(19)+in_buf[709]*(3)+in_buf[710]*(-10)+in_buf[711]*(-7)+in_buf[712]*(0)+in_buf[713]*(-6)+in_buf[714]*(8)+in_buf[715]*(5)+in_buf[716]*(-8)+in_buf[717]*(-1)+in_buf[718]*(1)+in_buf[719]*(-24)+in_buf[720]*(-23)+in_buf[721]*(-41)+in_buf[722]*(-17)+in_buf[723]*(-21)+in_buf[724]*(-29)+in_buf[725]*(-16)+in_buf[726]*(4)+in_buf[727]*(-2)+in_buf[728]*(3)+in_buf[729]*(1)+in_buf[730]*(0)+in_buf[731]*(-12)+in_buf[732]*(-41)+in_buf[733]*(-37)+in_buf[734]*(-15)+in_buf[735]*(14)+in_buf[736]*(4)+in_buf[737]*(6)+in_buf[738]*(-17)+in_buf[739]*(-8)+in_buf[740]*(-8)+in_buf[741]*(-3)+in_buf[742]*(-7)+in_buf[743]*(2)+in_buf[744]*(-13)+in_buf[745]*(-9)+in_buf[746]*(-7)+in_buf[747]*(-12)+in_buf[748]*(-7)+in_buf[749]*(-34)+in_buf[750]*(-38)+in_buf[751]*(-2)+in_buf[752]*(-23)+in_buf[753]*(11)+in_buf[754]*(-2)+in_buf[755]*(-1)+in_buf[756]*(0)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(0)+in_buf[760]*(35)+in_buf[761]*(21)+in_buf[762]*(13)+in_buf[763]*(3)+in_buf[764]*(5)+in_buf[765]*(23)+in_buf[766]*(7)+in_buf[767]*(0)+in_buf[768]*(1)+in_buf[769]*(41)+in_buf[770]*(-5)+in_buf[771]*(-10)+in_buf[772]*(18)+in_buf[773]*(39)+in_buf[774]*(22)+in_buf[775]*(-4)+in_buf[776]*(-10)+in_buf[777]*(-22)+in_buf[778]*(-21)+in_buf[779]*(-1)+in_buf[780]*(0)+in_buf[781]*(-2)+in_buf[782]*(-1)+in_buf[783]*(0);
assign in_buf_weight054=in_buf[0]*(4)+in_buf[1]*(0)+in_buf[2]*(3)+in_buf[3]*(0)+in_buf[4]*(1)+in_buf[5]*(-3)+in_buf[6]*(0)+in_buf[7]*(-2)+in_buf[8]*(-1)+in_buf[9]*(-2)+in_buf[10]*(0)+in_buf[11]*(0)+in_buf[12]*(-2)+in_buf[13]*(2)+in_buf[14]*(-1)+in_buf[15]*(-2)+in_buf[16]*(2)+in_buf[17]*(0)+in_buf[18]*(-3)+in_buf[19]*(0)+in_buf[20]*(-3)+in_buf[21]*(2)+in_buf[22]*(0)+in_buf[23]*(3)+in_buf[24]*(2)+in_buf[25]*(0)+in_buf[26]*(3)+in_buf[27]*(-2)+in_buf[28]*(-1)+in_buf[29]*(-1)+in_buf[30]*(4)+in_buf[31]*(1)+in_buf[32]*(0)+in_buf[33]*(8)+in_buf[34]*(5)+in_buf[35]*(8)+in_buf[36]*(13)+in_buf[37]*(9)+in_buf[38]*(1)+in_buf[39]*(14)+in_buf[40]*(24)+in_buf[41]*(15)+in_buf[42]*(-31)+in_buf[43]*(11)+in_buf[44]*(22)+in_buf[45]*(19)+in_buf[46]*(-2)+in_buf[47]*(-1)+in_buf[48]*(2)+in_buf[49]*(5)+in_buf[50]*(4)+in_buf[51]*(0)+in_buf[52]*(1)+in_buf[53]*(2)+in_buf[54]*(-1)+in_buf[55]*(-3)+in_buf[56]*(-1)+in_buf[57]*(2)+in_buf[58]*(5)+in_buf[59]*(28)+in_buf[60]*(36)+in_buf[61]*(7)+in_buf[62]*(7)+in_buf[63]*(15)+in_buf[64]*(2)+in_buf[65]*(24)+in_buf[66]*(35)+in_buf[67]*(31)+in_buf[68]*(27)+in_buf[69]*(-16)+in_buf[70]*(-24)+in_buf[71]*(-21)+in_buf[72]*(-1)+in_buf[73]*(-9)+in_buf[74]*(-30)+in_buf[75]*(-25)+in_buf[76]*(-51)+in_buf[77]*(-33)+in_buf[78]*(-30)+in_buf[79]*(12)+in_buf[80]*(5)+in_buf[81]*(4)+in_buf[82]*(2)+in_buf[83]*(-3)+in_buf[84]*(-3)+in_buf[85]*(2)+in_buf[86]*(-1)+in_buf[87]*(37)+in_buf[88]*(18)+in_buf[89]*(-7)+in_buf[90]*(-5)+in_buf[91]*(-17)+in_buf[92]*(0)+in_buf[93]*(-2)+in_buf[94]*(1)+in_buf[95]*(2)+in_buf[96]*(9)+in_buf[97]*(12)+in_buf[98]*(51)+in_buf[99]*(39)+in_buf[100]*(39)+in_buf[101]*(27)+in_buf[102]*(23)+in_buf[103]*(21)+in_buf[104]*(38)+in_buf[105]*(8)+in_buf[106]*(-22)+in_buf[107]*(-5)+in_buf[108]*(7)+in_buf[109]*(24)+in_buf[110]*(20)+in_buf[111]*(0)+in_buf[112]*(-1)+in_buf[113]*(4)+in_buf[114]*(23)+in_buf[115]*(13)+in_buf[116]*(18)+in_buf[117]*(5)+in_buf[118]*(1)+in_buf[119]*(-15)+in_buf[120]*(-28)+in_buf[121]*(-12)+in_buf[122]*(-16)+in_buf[123]*(13)+in_buf[124]*(17)+in_buf[125]*(19)+in_buf[126]*(13)+in_buf[127]*(22)+in_buf[128]*(20)+in_buf[129]*(27)+in_buf[130]*(21)+in_buf[131]*(8)+in_buf[132]*(10)+in_buf[133]*(3)+in_buf[134]*(6)+in_buf[135]*(-24)+in_buf[136]*(-31)+in_buf[137]*(-1)+in_buf[138]*(32)+in_buf[139]*(1)+in_buf[140]*(2)+in_buf[141]*(3)+in_buf[142]*(18)+in_buf[143]*(1)+in_buf[144]*(11)+in_buf[145]*(21)+in_buf[146]*(16)+in_buf[147]*(-13)+in_buf[148]*(-3)+in_buf[149]*(-16)+in_buf[150]*(-34)+in_buf[151]*(-25)+in_buf[152]*(-5)+in_buf[153]*(19)+in_buf[154]*(2)+in_buf[155]*(-2)+in_buf[156]*(8)+in_buf[157]*(-7)+in_buf[158]*(2)+in_buf[159]*(-11)+in_buf[160]*(-16)+in_buf[161]*(-7)+in_buf[162]*(9)+in_buf[163]*(-11)+in_buf[164]*(-33)+in_buf[165]*(-11)+in_buf[166]*(16)+in_buf[167]*(-14)+in_buf[168]*(-3)+in_buf[169]*(18)+in_buf[170]*(18)+in_buf[171]*(36)+in_buf[172]*(37)+in_buf[173]*(26)+in_buf[174]*(16)+in_buf[175]*(-10)+in_buf[176]*(-10)+in_buf[177]*(-27)+in_buf[178]*(-12)+in_buf[179]*(-11)+in_buf[180]*(-16)+in_buf[181]*(-10)+in_buf[182]*(-36)+in_buf[183]*(-38)+in_buf[184]*(-20)+in_buf[185]*(-3)+in_buf[186]*(5)+in_buf[187]*(0)+in_buf[188]*(-4)+in_buf[189]*(28)+in_buf[190]*(12)+in_buf[191]*(-1)+in_buf[192]*(1)+in_buf[193]*(-37)+in_buf[194]*(17)+in_buf[195]*(15)+in_buf[196]*(-2)+in_buf[197]*(39)+in_buf[198]*(19)+in_buf[199]*(54)+in_buf[200]*(17)+in_buf[201]*(0)+in_buf[202]*(6)+in_buf[203]*(3)+in_buf[204]*(-9)+in_buf[205]*(1)+in_buf[206]*(0)+in_buf[207]*(-6)+in_buf[208]*(-3)+in_buf[209]*(-19)+in_buf[210]*(-26)+in_buf[211]*(-20)+in_buf[212]*(-12)+in_buf[213]*(5)+in_buf[214]*(24)+in_buf[215]*(13)+in_buf[216]*(16)+in_buf[217]*(18)+in_buf[218]*(17)+in_buf[219]*(26)+in_buf[220]*(12)+in_buf[221]*(-14)+in_buf[222]*(-9)+in_buf[223]*(35)+in_buf[224]*(30)+in_buf[225]*(31)+in_buf[226]*(20)+in_buf[227]*(32)+in_buf[228]*(13)+in_buf[229]*(18)+in_buf[230]*(8)+in_buf[231]*(18)+in_buf[232]*(19)+in_buf[233]*(10)+in_buf[234]*(9)+in_buf[235]*(1)+in_buf[236]*(17)+in_buf[237]*(-5)+in_buf[238]*(10)+in_buf[239]*(15)+in_buf[240]*(12)+in_buf[241]*(20)+in_buf[242]*(27)+in_buf[243]*(18)+in_buf[244]*(18)+in_buf[245]*(13)+in_buf[246]*(35)+in_buf[247]*(32)+in_buf[248]*(6)+in_buf[249]*(-29)+in_buf[250]*(-29)+in_buf[251]*(12)+in_buf[252]*(10)+in_buf[253]*(36)+in_buf[254]*(2)+in_buf[255]*(13)+in_buf[256]*(7)+in_buf[257]*(18)+in_buf[258]*(15)+in_buf[259]*(19)+in_buf[260]*(11)+in_buf[261]*(8)+in_buf[262]*(14)+in_buf[263]*(4)+in_buf[264]*(27)+in_buf[265]*(20)+in_buf[266]*(24)+in_buf[267]*(20)+in_buf[268]*(26)+in_buf[269]*(31)+in_buf[270]*(21)+in_buf[271]*(26)+in_buf[272]*(23)+in_buf[273]*(8)+in_buf[274]*(29)+in_buf[275]*(33)+in_buf[276]*(11)+in_buf[277]*(-3)+in_buf[278]*(-24)+in_buf[279]*(7)+in_buf[280]*(19)+in_buf[281]*(24)+in_buf[282]*(39)+in_buf[283]*(-1)+in_buf[284]*(-9)+in_buf[285]*(-17)+in_buf[286]*(10)+in_buf[287]*(8)+in_buf[288]*(2)+in_buf[289]*(9)+in_buf[290]*(9)+in_buf[291]*(10)+in_buf[292]*(0)+in_buf[293]*(26)+in_buf[294]*(22)+in_buf[295]*(23)+in_buf[296]*(33)+in_buf[297]*(15)+in_buf[298]*(15)+in_buf[299]*(10)+in_buf[300]*(24)+in_buf[301]*(8)+in_buf[302]*(21)+in_buf[303]*(-5)+in_buf[304]*(5)+in_buf[305]*(-3)+in_buf[306]*(-1)+in_buf[307]*(-14)+in_buf[308]*(15)+in_buf[309]*(36)+in_buf[310]*(35)+in_buf[311]*(0)+in_buf[312]*(-29)+in_buf[313]*(-40)+in_buf[314]*(-5)+in_buf[315]*(12)+in_buf[316]*(0)+in_buf[317]*(0)+in_buf[318]*(9)+in_buf[319]*(6)+in_buf[320]*(4)+in_buf[321]*(14)+in_buf[322]*(14)+in_buf[323]*(4)+in_buf[324]*(-10)+in_buf[325]*(-6)+in_buf[326]*(13)+in_buf[327]*(0)+in_buf[328]*(9)+in_buf[329]*(-5)+in_buf[330]*(-9)+in_buf[331]*(-16)+in_buf[332]*(-15)+in_buf[333]*(-32)+in_buf[334]*(-2)+in_buf[335]*(6)+in_buf[336]*(24)+in_buf[337]*(14)+in_buf[338]*(6)+in_buf[339]*(-10)+in_buf[340]*(-41)+in_buf[341]*(-33)+in_buf[342]*(-7)+in_buf[343]*(8)+in_buf[344]*(4)+in_buf[345]*(1)+in_buf[346]*(3)+in_buf[347]*(-1)+in_buf[348]*(-2)+in_buf[349]*(-13)+in_buf[350]*(-5)+in_buf[351]*(-15)+in_buf[352]*(-23)+in_buf[353]*(-11)+in_buf[354]*(1)+in_buf[355]*(-1)+in_buf[356]*(0)+in_buf[357]*(-10)+in_buf[358]*(-1)+in_buf[359]*(-12)+in_buf[360]*(-18)+in_buf[361]*(-34)+in_buf[362]*(-42)+in_buf[363]*(-22)+in_buf[364]*(2)+in_buf[365]*(9)+in_buf[366]*(33)+in_buf[367]*(3)+in_buf[368]*(-25)+in_buf[369]*(-5)+in_buf[370]*(5)+in_buf[371]*(4)+in_buf[372]*(8)+in_buf[373]*(0)+in_buf[374]*(-6)+in_buf[375]*(-21)+in_buf[376]*(-22)+in_buf[377]*(-29)+in_buf[378]*(-15)+in_buf[379]*(-31)+in_buf[380]*(-15)+in_buf[381]*(-7)+in_buf[382]*(3)+in_buf[383]*(4)+in_buf[384]*(-1)+in_buf[385]*(3)+in_buf[386]*(-1)+in_buf[387]*(-3)+in_buf[388]*(1)+in_buf[389]*(-14)+in_buf[390]*(-50)+in_buf[391]*(-24)+in_buf[392]*(14)+in_buf[393]*(14)+in_buf[394]*(29)+in_buf[395]*(4)+in_buf[396]*(-14)+in_buf[397]*(3)+in_buf[398]*(5)+in_buf[399]*(7)+in_buf[400]*(3)+in_buf[401]*(0)+in_buf[402]*(-15)+in_buf[403]*(-19)+in_buf[404]*(-22)+in_buf[405]*(-27)+in_buf[406]*(-15)+in_buf[407]*(-9)+in_buf[408]*(-19)+in_buf[409]*(-1)+in_buf[410]*(9)+in_buf[411]*(5)+in_buf[412]*(2)+in_buf[413]*(2)+in_buf[414]*(-5)+in_buf[415]*(13)+in_buf[416]*(30)+in_buf[417]*(-12)+in_buf[418]*(-30)+in_buf[419]*(-16)+in_buf[420]*(8)+in_buf[421]*(6)+in_buf[422]*(10)+in_buf[423]*(-18)+in_buf[424]*(-10)+in_buf[425]*(11)+in_buf[426]*(17)+in_buf[427]*(11)+in_buf[428]*(-12)+in_buf[429]*(-20)+in_buf[430]*(-29)+in_buf[431]*(-43)+in_buf[432]*(-19)+in_buf[433]*(-36)+in_buf[434]*(-14)+in_buf[435]*(-5)+in_buf[436]*(-22)+in_buf[437]*(-2)+in_buf[438]*(3)+in_buf[439]*(-3)+in_buf[440]*(4)+in_buf[441]*(10)+in_buf[442]*(7)+in_buf[443]*(17)+in_buf[444]*(37)+in_buf[445]*(-9)+in_buf[446]*(-15)+in_buf[447]*(-14)+in_buf[448]*(3)+in_buf[449]*(7)+in_buf[450]*(11)+in_buf[451]*(-15)+in_buf[452]*(3)+in_buf[453]*(12)+in_buf[454]*(2)+in_buf[455]*(6)+in_buf[456]*(8)+in_buf[457]*(-10)+in_buf[458]*(-30)+in_buf[459]*(-32)+in_buf[460]*(-21)+in_buf[461]*(-16)+in_buf[462]*(-10)+in_buf[463]*(-6)+in_buf[464]*(-14)+in_buf[465]*(7)+in_buf[466]*(4)+in_buf[467]*(-5)+in_buf[468]*(6)+in_buf[469]*(-13)+in_buf[470]*(-17)+in_buf[471]*(-8)+in_buf[472]*(9)+in_buf[473]*(-42)+in_buf[474]*(-23)+in_buf[475]*(5)+in_buf[476]*(2)+in_buf[477]*(13)+in_buf[478]*(-21)+in_buf[479]*(-7)+in_buf[480]*(9)+in_buf[481]*(0)+in_buf[482]*(0)+in_buf[483]*(15)+in_buf[484]*(15)+in_buf[485]*(9)+in_buf[486]*(-7)+in_buf[487]*(-3)+in_buf[488]*(-11)+in_buf[489]*(-2)+in_buf[490]*(-4)+in_buf[491]*(0)+in_buf[492]*(-2)+in_buf[493]*(17)+in_buf[494]*(3)+in_buf[495]*(7)+in_buf[496]*(-6)+in_buf[497]*(-19)+in_buf[498]*(-12)+in_buf[499]*(2)+in_buf[500]*(6)+in_buf[501]*(-2)+in_buf[502]*(-29)+in_buf[503]*(18)+in_buf[504]*(31)+in_buf[505]*(10)+in_buf[506]*(-6)+in_buf[507]*(-17)+in_buf[508]*(-11)+in_buf[509]*(4)+in_buf[510]*(3)+in_buf[511]*(16)+in_buf[512]*(34)+in_buf[513]*(20)+in_buf[514]*(8)+in_buf[515]*(9)+in_buf[516]*(-9)+in_buf[517]*(-6)+in_buf[518]*(0)+in_buf[519]*(11)+in_buf[520]*(10)+in_buf[521]*(19)+in_buf[522]*(16)+in_buf[523]*(-5)+in_buf[524]*(4)+in_buf[525]*(-3)+in_buf[526]*(7)+in_buf[527]*(-1)+in_buf[528]*(-4)+in_buf[529]*(3)+in_buf[530]*(-13)+in_buf[531]*(-8)+in_buf[532]*(1)+in_buf[533]*(47)+in_buf[534]*(45)+in_buf[535]*(-23)+in_buf[536]*(4)+in_buf[537]*(5)+in_buf[538]*(0)+in_buf[539]*(1)+in_buf[540]*(27)+in_buf[541]*(18)+in_buf[542]*(3)+in_buf[543]*(-5)+in_buf[544]*(-4)+in_buf[545]*(2)+in_buf[546]*(8)+in_buf[547]*(-7)+in_buf[548]*(-8)+in_buf[549]*(3)+in_buf[550]*(-9)+in_buf[551]*(-11)+in_buf[552]*(-8)+in_buf[553]*(-20)+in_buf[554]*(-11)+in_buf[555]*(-23)+in_buf[556]*(-15)+in_buf[557]*(-19)+in_buf[558]*(-17)+in_buf[559]*(-6)+in_buf[560]*(0)+in_buf[561]*(26)+in_buf[562]*(6)+in_buf[563]*(-17)+in_buf[564]*(6)+in_buf[565]*(0)+in_buf[566]*(-12)+in_buf[567]*(-4)+in_buf[568]*(13)+in_buf[569]*(8)+in_buf[570]*(2)+in_buf[571]*(-1)+in_buf[572]*(10)+in_buf[573]*(17)+in_buf[574]*(14)+in_buf[575]*(-2)+in_buf[576]*(-16)+in_buf[577]*(-9)+in_buf[578]*(-30)+in_buf[579]*(-28)+in_buf[580]*(-29)+in_buf[581]*(-47)+in_buf[582]*(-37)+in_buf[583]*(-33)+in_buf[584]*(-24)+in_buf[585]*(-9)+in_buf[586]*(-10)+in_buf[587]*(4)+in_buf[588]*(-17)+in_buf[589]*(4)+in_buf[590]*(-8)+in_buf[591]*(-25)+in_buf[592]*(-9)+in_buf[593]*(-17)+in_buf[594]*(-21)+in_buf[595]*(-11)+in_buf[596]*(-11)+in_buf[597]*(-5)+in_buf[598]*(0)+in_buf[599]*(0)+in_buf[600]*(14)+in_buf[601]*(12)+in_buf[602]*(4)+in_buf[603]*(-4)+in_buf[604]*(-11)+in_buf[605]*(-7)+in_buf[606]*(-23)+in_buf[607]*(-33)+in_buf[608]*(-60)+in_buf[609]*(-40)+in_buf[610]*(-40)+in_buf[611]*(-43)+in_buf[612]*(-21)+in_buf[613]*(-21)+in_buf[614]*(29)+in_buf[615]*(7)+in_buf[616]*(-10)+in_buf[617]*(7)+in_buf[618]*(7)+in_buf[619]*(-15)+in_buf[620]*(-11)+in_buf[621]*(-16)+in_buf[622]*(-9)+in_buf[623]*(1)+in_buf[624]*(-6)+in_buf[625]*(1)+in_buf[626]*(-6)+in_buf[627]*(-11)+in_buf[628]*(9)+in_buf[629]*(11)+in_buf[630]*(8)+in_buf[631]*(-5)+in_buf[632]*(3)+in_buf[633]*(0)+in_buf[634]*(-33)+in_buf[635]*(-59)+in_buf[636]*(-47)+in_buf[637]*(-44)+in_buf[638]*(-46)+in_buf[639]*(-51)+in_buf[640]*(-44)+in_buf[641]*(-1)+in_buf[642]*(25)+in_buf[643]*(3)+in_buf[644]*(0)+in_buf[645]*(0)+in_buf[646]*(24)+in_buf[647]*(7)+in_buf[648]*(7)+in_buf[649]*(11)+in_buf[650]*(6)+in_buf[651]*(7)+in_buf[652]*(-18)+in_buf[653]*(-11)+in_buf[654]*(7)+in_buf[655]*(22)+in_buf[656]*(14)+in_buf[657]*(6)+in_buf[658]*(0)+in_buf[659]*(-11)+in_buf[660]*(0)+in_buf[661]*(-2)+in_buf[662]*(-33)+in_buf[663]*(-70)+in_buf[664]*(-43)+in_buf[665]*(-29)+in_buf[666]*(-21)+in_buf[667]*(-17)+in_buf[668]*(-30)+in_buf[669]*(-3)+in_buf[670]*(-8)+in_buf[671]*(0)+in_buf[672]*(4)+in_buf[673]*(1)+in_buf[674]*(14)+in_buf[675]*(38)+in_buf[676]*(53)+in_buf[677]*(37)+in_buf[678]*(5)+in_buf[679]*(-4)+in_buf[680]*(-14)+in_buf[681]*(-12)+in_buf[682]*(3)+in_buf[683]*(15)+in_buf[684]*(13)+in_buf[685]*(8)+in_buf[686]*(1)+in_buf[687]*(0)+in_buf[688]*(0)+in_buf[689]*(-16)+in_buf[690]*(-48)+in_buf[691]*(-48)+in_buf[692]*(-18)+in_buf[693]*(-14)+in_buf[694]*(-31)+in_buf[695]*(-26)+in_buf[696]*(-12)+in_buf[697]*(-19)+in_buf[698]*(-3)+in_buf[699]*(2)+in_buf[700]*(3)+in_buf[701]*(0)+in_buf[702]*(-33)+in_buf[703]*(27)+in_buf[704]*(28)+in_buf[705]*(12)+in_buf[706]*(13)+in_buf[707]*(28)+in_buf[708]*(8)+in_buf[709]*(2)+in_buf[710]*(15)+in_buf[711]*(16)+in_buf[712]*(11)+in_buf[713]*(-6)+in_buf[714]*(-6)+in_buf[715]*(5)+in_buf[716]*(19)+in_buf[717]*(-8)+in_buf[718]*(-17)+in_buf[719]*(-13)+in_buf[720]*(3)+in_buf[721]*(10)+in_buf[722]*(3)+in_buf[723]*(3)+in_buf[724]*(9)+in_buf[725]*(-3)+in_buf[726]*(-3)+in_buf[727]*(3)+in_buf[728]*(1)+in_buf[729]*(0)+in_buf[730]*(2)+in_buf[731]*(1)+in_buf[732]*(-39)+in_buf[733]*(-36)+in_buf[734]*(-21)+in_buf[735]*(12)+in_buf[736]*(10)+in_buf[737]*(24)+in_buf[738]*(9)+in_buf[739]*(11)+in_buf[740]*(8)+in_buf[741]*(35)+in_buf[742]*(14)+in_buf[743]*(5)+in_buf[744]*(11)+in_buf[745]*(-5)+in_buf[746]*(4)+in_buf[747]*(26)+in_buf[748]*(23)+in_buf[749]*(20)+in_buf[750]*(4)+in_buf[751]*(0)+in_buf[752]*(-28)+in_buf[753]*(12)+in_buf[754]*(2)+in_buf[755]*(3)+in_buf[756]*(-2)+in_buf[757]*(2)+in_buf[758]*(2)+in_buf[759]*(4)+in_buf[760]*(26)+in_buf[761]*(45)+in_buf[762]*(23)+in_buf[763]*(4)+in_buf[764]*(10)+in_buf[765]*(22)+in_buf[766]*(28)+in_buf[767]*(22)+in_buf[768]*(11)+in_buf[769]*(51)+in_buf[770]*(28)+in_buf[771]*(-8)+in_buf[772]*(7)+in_buf[773]*(44)+in_buf[774]*(25)+in_buf[775]*(3)+in_buf[776]*(8)+in_buf[777]*(11)+in_buf[778]*(0)+in_buf[779]*(24)+in_buf[780]*(0)+in_buf[781]*(1)+in_buf[782]*(-2)+in_buf[783]*(4);
assign in_buf_weight055=in_buf[0]*(1)+in_buf[1]*(0)+in_buf[2]*(0)+in_buf[3]*(4)+in_buf[4]*(0)+in_buf[5]*(4)+in_buf[6]*(0)+in_buf[7]*(0)+in_buf[8]*(1)+in_buf[9]*(0)+in_buf[10]*(2)+in_buf[11]*(2)+in_buf[12]*(12)+in_buf[13]*(9)+in_buf[14]*(7)+in_buf[15]*(2)+in_buf[16]*(0)+in_buf[17]*(3)+in_buf[18]*(2)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(4)+in_buf[22]*(-3)+in_buf[23]*(-2)+in_buf[24]*(0)+in_buf[25]*(3)+in_buf[26]*(-3)+in_buf[27]*(0)+in_buf[28]*(0)+in_buf[29]*(0)+in_buf[30]*(-3)+in_buf[31]*(3)+in_buf[32]*(5)+in_buf[33]*(0)+in_buf[34]*(-6)+in_buf[35]*(-11)+in_buf[36]*(-3)+in_buf[37]*(-5)+in_buf[38]*(-19)+in_buf[39]*(-4)+in_buf[40]*(-4)+in_buf[41]*(24)+in_buf[42]*(23)+in_buf[43]*(18)+in_buf[44]*(19)+in_buf[45]*(18)+in_buf[46]*(-1)+in_buf[47]*(-7)+in_buf[48]*(2)+in_buf[49]*(7)+in_buf[50]*(-12)+in_buf[51]*(-4)+in_buf[52]*(-1)+in_buf[53]*(3)+in_buf[54]*(0)+in_buf[55]*(4)+in_buf[56]*(-1)+in_buf[57]*(2)+in_buf[58]*(8)+in_buf[59]*(19)+in_buf[60]*(25)+in_buf[61]*(-5)+in_buf[62]*(-8)+in_buf[63]*(-20)+in_buf[64]*(-14)+in_buf[65]*(-42)+in_buf[66]*(-46)+in_buf[67]*(-18)+in_buf[68]*(2)+in_buf[69]*(-9)+in_buf[70]*(-2)+in_buf[71]*(-19)+in_buf[72]*(-1)+in_buf[73]*(-6)+in_buf[74]*(-1)+in_buf[75]*(-12)+in_buf[76]*(-11)+in_buf[77]*(-23)+in_buf[78]*(-15)+in_buf[79]*(9)+in_buf[80]*(-25)+in_buf[81]*(0)+in_buf[82]*(-2)+in_buf[83]*(1)+in_buf[84]*(-3)+in_buf[85]*(0)+in_buf[86]*(9)+in_buf[87]*(19)+in_buf[88]*(15)+in_buf[89]*(8)+in_buf[90]*(-7)+in_buf[91]*(0)+in_buf[92]*(16)+in_buf[93]*(-4)+in_buf[94]*(14)+in_buf[95]*(15)+in_buf[96]*(20)+in_buf[97]*(8)+in_buf[98]*(14)+in_buf[99]*(15)+in_buf[100]*(15)+in_buf[101]*(8)+in_buf[102]*(9)+in_buf[103]*(13)+in_buf[104]*(53)+in_buf[105]*(29)+in_buf[106]*(-14)+in_buf[107]*(10)+in_buf[108]*(23)+in_buf[109]*(10)+in_buf[110]*(0)+in_buf[111]*(-2)+in_buf[112]*(-3)+in_buf[113]*(5)+in_buf[114]*(11)+in_buf[115]*(16)+in_buf[116]*(4)+in_buf[117]*(0)+in_buf[118]*(-11)+in_buf[119]*(12)+in_buf[120]*(10)+in_buf[121]*(7)+in_buf[122]*(18)+in_buf[123]*(21)+in_buf[124]*(20)+in_buf[125]*(8)+in_buf[126]*(12)+in_buf[127]*(16)+in_buf[128]*(10)+in_buf[129]*(-1)+in_buf[130]*(1)+in_buf[131]*(7)+in_buf[132]*(12)+in_buf[133]*(24)+in_buf[134]*(-5)+in_buf[135]*(-31)+in_buf[136]*(5)+in_buf[137]*(12)+in_buf[138]*(13)+in_buf[139]*(15)+in_buf[140]*(0)+in_buf[141]*(-2)+in_buf[142]*(-2)+in_buf[143]*(7)+in_buf[144]*(-17)+in_buf[145]*(0)+in_buf[146]*(3)+in_buf[147]*(27)+in_buf[148]*(9)+in_buf[149]*(17)+in_buf[150]*(3)+in_buf[151]*(12)+in_buf[152]*(7)+in_buf[153]*(9)+in_buf[154]*(6)+in_buf[155]*(3)+in_buf[156]*(8)+in_buf[157]*(13)+in_buf[158]*(6)+in_buf[159]*(-3)+in_buf[160]*(-5)+in_buf[161]*(-11)+in_buf[162]*(-40)+in_buf[163]*(-52)+in_buf[164]*(-35)+in_buf[165]*(-9)+in_buf[166]*(35)+in_buf[167]*(20)+in_buf[168]*(3)+in_buf[169]*(-5)+in_buf[170]*(10)+in_buf[171]*(7)+in_buf[172]*(5)+in_buf[173]*(4)+in_buf[174]*(9)+in_buf[175]*(9)+in_buf[176]*(16)+in_buf[177]*(9)+in_buf[178]*(3)+in_buf[179]*(4)+in_buf[180]*(-4)+in_buf[181]*(0)+in_buf[182]*(4)+in_buf[183]*(9)+in_buf[184]*(7)+in_buf[185]*(16)+in_buf[186]*(12)+in_buf[187]*(4)+in_buf[188]*(9)+in_buf[189]*(13)+in_buf[190]*(-12)+in_buf[191]*(-26)+in_buf[192]*(-11)+in_buf[193]*(13)+in_buf[194]*(23)+in_buf[195]*(3)+in_buf[196]*(-2)+in_buf[197]*(18)+in_buf[198]*(3)+in_buf[199]*(18)+in_buf[200]*(-6)+in_buf[201]*(-20)+in_buf[202]*(0)+in_buf[203]*(13)+in_buf[204]*(0)+in_buf[205]*(8)+in_buf[206]*(8)+in_buf[207]*(-7)+in_buf[208]*(-5)+in_buf[209]*(-9)+in_buf[210]*(-14)+in_buf[211]*(4)+in_buf[212]*(-1)+in_buf[213]*(0)+in_buf[214]*(7)+in_buf[215]*(0)+in_buf[216]*(2)+in_buf[217]*(-4)+in_buf[218]*(-5)+in_buf[219]*(2)+in_buf[220]*(10)+in_buf[221]*(25)+in_buf[222]*(22)+in_buf[223]*(11)+in_buf[224]*(-24)+in_buf[225]*(26)+in_buf[226]*(12)+in_buf[227]*(18)+in_buf[228]*(-9)+in_buf[229]*(-10)+in_buf[230]*(-10)+in_buf[231]*(1)+in_buf[232]*(1)+in_buf[233]*(-6)+in_buf[234]*(6)+in_buf[235]*(0)+in_buf[236]*(7)+in_buf[237]*(-3)+in_buf[238]*(-1)+in_buf[239]*(0)+in_buf[240]*(-5)+in_buf[241]*(-13)+in_buf[242]*(7)+in_buf[243]*(6)+in_buf[244]*(9)+in_buf[245]*(17)+in_buf[246]*(19)+in_buf[247]*(11)+in_buf[248]*(47)+in_buf[249]*(34)+in_buf[250]*(-7)+in_buf[251]*(32)+in_buf[252]*(17)+in_buf[253]*(30)+in_buf[254]*(13)+in_buf[255]*(7)+in_buf[256]*(13)+in_buf[257]*(1)+in_buf[258]*(1)+in_buf[259]*(-10)+in_buf[260]*(-8)+in_buf[261]*(6)+in_buf[262]*(11)+in_buf[263]*(7)+in_buf[264]*(4)+in_buf[265]*(13)+in_buf[266]*(15)+in_buf[267]*(-7)+in_buf[268]*(-8)+in_buf[269]*(5)+in_buf[270]*(6)+in_buf[271]*(13)+in_buf[272]*(32)+in_buf[273]*(25)+in_buf[274]*(29)+in_buf[275]*(22)+in_buf[276]*(29)+in_buf[277]*(60)+in_buf[278]*(24)+in_buf[279]*(26)+in_buf[280]*(17)+in_buf[281]*(14)+in_buf[282]*(18)+in_buf[283]*(13)+in_buf[284]*(24)+in_buf[285]*(-6)+in_buf[286]*(0)+in_buf[287]*(-12)+in_buf[288]*(-14)+in_buf[289]*(12)+in_buf[290]*(6)+in_buf[291]*(6)+in_buf[292]*(6)+in_buf[293]*(16)+in_buf[294]*(26)+in_buf[295]*(4)+in_buf[296]*(4)+in_buf[297]*(-1)+in_buf[298]*(6)+in_buf[299]*(16)+in_buf[300]*(43)+in_buf[301]*(19)+in_buf[302]*(24)+in_buf[303]*(18)+in_buf[304]*(10)+in_buf[305]*(55)+in_buf[306]*(41)+in_buf[307]*(26)+in_buf[308]*(22)+in_buf[309]*(4)+in_buf[310]*(39)+in_buf[311]*(38)+in_buf[312]*(24)+in_buf[313]*(-8)+in_buf[314]*(-15)+in_buf[315]*(-20)+in_buf[316]*(1)+in_buf[317]*(6)+in_buf[318]*(-3)+in_buf[319]*(7)+in_buf[320]*(23)+in_buf[321]*(31)+in_buf[322]*(31)+in_buf[323]*(17)+in_buf[324]*(8)+in_buf[325]*(14)+in_buf[326]*(21)+in_buf[327]*(17)+in_buf[328]*(32)+in_buf[329]*(10)+in_buf[330]*(10)+in_buf[331]*(-1)+in_buf[332]*(-3)+in_buf[333]*(37)+in_buf[334]*(12)+in_buf[335]*(-8)+in_buf[336]*(22)+in_buf[337]*(10)+in_buf[338]*(25)+in_buf[339]*(40)+in_buf[340]*(25)+in_buf[341]*(4)+in_buf[342]*(-18)+in_buf[343]*(-5)+in_buf[344]*(-1)+in_buf[345]*(-6)+in_buf[346]*(-10)+in_buf[347]*(10)+in_buf[348]*(7)+in_buf[349]*(22)+in_buf[350]*(26)+in_buf[351]*(28)+in_buf[352]*(17)+in_buf[353]*(16)+in_buf[354]*(18)+in_buf[355]*(15)+in_buf[356]*(8)+in_buf[357]*(-12)+in_buf[358]*(-21)+in_buf[359]*(-34)+in_buf[360]*(-63)+in_buf[361]*(-22)+in_buf[362]*(11)+in_buf[363]*(-2)+in_buf[364]*(-21)+in_buf[365]*(0)+in_buf[366]*(30)+in_buf[367]*(29)+in_buf[368]*(30)+in_buf[369]*(21)+in_buf[370]*(-1)+in_buf[371]*(-9)+in_buf[372]*(-12)+in_buf[373]*(-15)+in_buf[374]*(-15)+in_buf[375]*(-9)+in_buf[376]*(-15)+in_buf[377]*(7)+in_buf[378]*(11)+in_buf[379]*(19)+in_buf[380]*(18)+in_buf[381]*(-2)+in_buf[382]*(5)+in_buf[383]*(0)+in_buf[384]*(4)+in_buf[385]*(-8)+in_buf[386]*(-35)+in_buf[387]*(-52)+in_buf[388]*(-58)+in_buf[389]*(-34)+in_buf[390]*(-8)+in_buf[391]*(-9)+in_buf[392]*(0)+in_buf[393]*(0)+in_buf[394]*(9)+in_buf[395]*(26)+in_buf[396]*(21)+in_buf[397]*(6)+in_buf[398]*(-9)+in_buf[399]*(-20)+in_buf[400]*(-16)+in_buf[401]*(-21)+in_buf[402]*(-15)+in_buf[403]*(-25)+in_buf[404]*(-15)+in_buf[405]*(-10)+in_buf[406]*(5)+in_buf[407]*(13)+in_buf[408]*(4)+in_buf[409]*(1)+in_buf[410]*(7)+in_buf[411]*(18)+in_buf[412]*(-1)+in_buf[413]*(-5)+in_buf[414]*(-28)+in_buf[415]*(2)+in_buf[416]*(-20)+in_buf[417]*(-31)+in_buf[418]*(-25)+in_buf[419]*(-8)+in_buf[420]*(10)+in_buf[421]*(2)+in_buf[422]*(-3)+in_buf[423]*(5)+in_buf[424]*(15)+in_buf[425]*(7)+in_buf[426]*(9)+in_buf[427]*(-1)+in_buf[428]*(-13)+in_buf[429]*(-25)+in_buf[430]*(-19)+in_buf[431]*(-22)+in_buf[432]*(-20)+in_buf[433]*(-13)+in_buf[434]*(-3)+in_buf[435]*(3)+in_buf[436]*(-6)+in_buf[437]*(6)+in_buf[438]*(18)+in_buf[439]*(25)+in_buf[440]*(24)+in_buf[441]*(-3)+in_buf[442]*(8)+in_buf[443]*(11)+in_buf[444]*(-32)+in_buf[445]*(-32)+in_buf[446]*(-13)+in_buf[447]*(-6)+in_buf[448]*(2)+in_buf[449]*(3)+in_buf[450]*(5)+in_buf[451]*(4)+in_buf[452]*(19)+in_buf[453]*(15)+in_buf[454]*(9)+in_buf[455]*(5)+in_buf[456]*(-12)+in_buf[457]*(-21)+in_buf[458]*(-24)+in_buf[459]*(-32)+in_buf[460]*(-17)+in_buf[461]*(-15)+in_buf[462]*(-15)+in_buf[463]*(-12)+in_buf[464]*(-14)+in_buf[465]*(10)+in_buf[466]*(17)+in_buf[467]*(9)+in_buf[468]*(17)+in_buf[469]*(-7)+in_buf[470]*(-14)+in_buf[471]*(-6)+in_buf[472]*(-24)+in_buf[473]*(-56)+in_buf[474]*(-25)+in_buf[475]*(-8)+in_buf[476]*(-1)+in_buf[477]*(13)+in_buf[478]*(-22)+in_buf[479]*(10)+in_buf[480]*(22)+in_buf[481]*(12)+in_buf[482]*(12)+in_buf[483]*(5)+in_buf[484]*(-9)+in_buf[485]*(-11)+in_buf[486]*(-18)+in_buf[487]*(-7)+in_buf[488]*(-13)+in_buf[489]*(-16)+in_buf[490]*(-22)+in_buf[491]*(-7)+in_buf[492]*(-13)+in_buf[493]*(5)+in_buf[494]*(9)+in_buf[495]*(5)+in_buf[496]*(1)+in_buf[497]*(-13)+in_buf[498]*(-18)+in_buf[499]*(-21)+in_buf[500]*(-28)+in_buf[501]*(-44)+in_buf[502]*(-16)+in_buf[503]*(11)+in_buf[504]*(32)+in_buf[505]*(8)+in_buf[506]*(-5)+in_buf[507]*(-9)+in_buf[508]*(10)+in_buf[509]*(12)+in_buf[510]*(12)+in_buf[511]*(9)+in_buf[512]*(-1)+in_buf[513]*(5)+in_buf[514]*(6)+in_buf[515]*(10)+in_buf[516]*(-7)+in_buf[517]*(-16)+in_buf[518]*(-20)+in_buf[519]*(-1)+in_buf[520]*(-1)+in_buf[521]*(10)+in_buf[522]*(19)+in_buf[523]*(12)+in_buf[524]*(10)+in_buf[525]*(-4)+in_buf[526]*(-27)+in_buf[527]*(-40)+in_buf[528]*(-53)+in_buf[529]*(-21)+in_buf[530]*(-3)+in_buf[531]*(-21)+in_buf[532]*(-19)+in_buf[533]*(32)+in_buf[534]*(12)+in_buf[535]*(-18)+in_buf[536]*(4)+in_buf[537]*(13)+in_buf[538]*(7)+in_buf[539]*(-5)+in_buf[540]*(0)+in_buf[541]*(-3)+in_buf[542]*(0)+in_buf[543]*(-4)+in_buf[544]*(-9)+in_buf[545]*(-19)+in_buf[546]*(-10)+in_buf[547]*(-5)+in_buf[548]*(4)+in_buf[549]*(10)+in_buf[550]*(10)+in_buf[551]*(4)+in_buf[552]*(0)+in_buf[553]*(-16)+in_buf[554]*(-39)+in_buf[555]*(-45)+in_buf[556]*(-32)+in_buf[557]*(-14)+in_buf[558]*(-9)+in_buf[559]*(-21)+in_buf[560]*(3)+in_buf[561]*(23)+in_buf[562]*(-24)+in_buf[563]*(-35)+in_buf[564]*(-3)+in_buf[565]*(-5)+in_buf[566]*(-9)+in_buf[567]*(-10)+in_buf[568]*(12)+in_buf[569]*(-1)+in_buf[570]*(-3)+in_buf[571]*(-15)+in_buf[572]*(-15)+in_buf[573]*(-4)+in_buf[574]*(-5)+in_buf[575]*(0)+in_buf[576]*(-4)+in_buf[577]*(0)+in_buf[578]*(-4)+in_buf[579]*(-2)+in_buf[580]*(-5)+in_buf[581]*(-21)+in_buf[582]*(-35)+in_buf[583]*(-46)+in_buf[584]*(-35)+in_buf[585]*(-25)+in_buf[586]*(-3)+in_buf[587]*(0)+in_buf[588]*(-28)+in_buf[589]*(-2)+in_buf[590]*(-23)+in_buf[591]*(-41)+in_buf[592]*(-15)+in_buf[593]*(-30)+in_buf[594]*(-11)+in_buf[595]*(-1)+in_buf[596]*(4)+in_buf[597]*(-8)+in_buf[598]*(-11)+in_buf[599]*(-1)+in_buf[600]*(-4)+in_buf[601]*(-7)+in_buf[602]*(-13)+in_buf[603]*(-4)+in_buf[604]*(-1)+in_buf[605]*(0)+in_buf[606]*(-12)+in_buf[607]*(-4)+in_buf[608]*(-5)+in_buf[609]*(-12)+in_buf[610]*(-41)+in_buf[611]*(-58)+in_buf[612]*(-31)+in_buf[613]*(-17)+in_buf[614]*(-23)+in_buf[615]*(2)+in_buf[616]*(-28)+in_buf[617]*(4)+in_buf[618]*(-20)+in_buf[619]*(-15)+in_buf[620]*(-3)+in_buf[621]*(-27)+in_buf[622]*(-15)+in_buf[623]*(-2)+in_buf[624]*(-7)+in_buf[625]*(-9)+in_buf[626]*(-12)+in_buf[627]*(-4)+in_buf[628]*(-6)+in_buf[629]*(-18)+in_buf[630]*(-2)+in_buf[631]*(1)+in_buf[632]*(0)+in_buf[633]*(-1)+in_buf[634]*(-21)+in_buf[635]*(-15)+in_buf[636]*(-33)+in_buf[637]*(-33)+in_buf[638]*(-36)+in_buf[639]*(-44)+in_buf[640]*(-37)+in_buf[641]*(-21)+in_buf[642]*(-34)+in_buf[643]*(-1)+in_buf[644]*(-3)+in_buf[645]*(-1)+in_buf[646]*(-14)+in_buf[647]*(19)+in_buf[648]*(26)+in_buf[649]*(-6)+in_buf[650]*(-26)+in_buf[651]*(-14)+in_buf[652]*(-11)+in_buf[653]*(-13)+in_buf[654]*(2)+in_buf[655]*(3)+in_buf[656]*(-9)+in_buf[657]*(-16)+in_buf[658]*(-5)+in_buf[659]*(-7)+in_buf[660]*(-1)+in_buf[661]*(-11)+in_buf[662]*(-19)+in_buf[663]*(-29)+in_buf[664]*(-38)+in_buf[665]*(-32)+in_buf[666]*(-37)+in_buf[667]*(-30)+in_buf[668]*(-21)+in_buf[669]*(-21)+in_buf[670]*(-35)+in_buf[671]*(-1)+in_buf[672]*(-2)+in_buf[673]*(-1)+in_buf[674]*(14)+in_buf[675]*(33)+in_buf[676]*(25)+in_buf[677]*(21)+in_buf[678]*(10)+in_buf[679]*(10)+in_buf[680]*(3)+in_buf[681]*(-13)+in_buf[682]*(2)+in_buf[683]*(-2)+in_buf[684]*(4)+in_buf[685]*(22)+in_buf[686]*(8)+in_buf[687]*(21)+in_buf[688]*(13)+in_buf[689]*(-6)+in_buf[690]*(-25)+in_buf[691]*(-13)+in_buf[692]*(-11)+in_buf[693]*(-44)+in_buf[694]*(-28)+in_buf[695]*(-29)+in_buf[696]*(-26)+in_buf[697]*(-21)+in_buf[698]*(-13)+in_buf[699]*(-1)+in_buf[700]*(0)+in_buf[701]*(3)+in_buf[702]*(31)+in_buf[703]*(7)+in_buf[704]*(9)+in_buf[705]*(11)+in_buf[706]*(8)+in_buf[707]*(20)+in_buf[708]*(11)+in_buf[709]*(14)+in_buf[710]*(16)+in_buf[711]*(22)+in_buf[712]*(35)+in_buf[713]*(38)+in_buf[714]*(5)+in_buf[715]*(25)+in_buf[716]*(29)+in_buf[717]*(3)+in_buf[718]*(-4)+in_buf[719]*(34)+in_buf[720]*(19)+in_buf[721]*(5)+in_buf[722]*(-9)+in_buf[723]*(-18)+in_buf[724]*(-1)+in_buf[725]*(11)+in_buf[726]*(0)+in_buf[727]*(-1)+in_buf[728]*(-1)+in_buf[729]*(-2)+in_buf[730]*(-3)+in_buf[731]*(22)+in_buf[732]*(-24)+in_buf[733]*(-17)+in_buf[734]*(-2)+in_buf[735]*(25)+in_buf[736]*(42)+in_buf[737]*(56)+in_buf[738]*(36)+in_buf[739]*(39)+in_buf[740]*(34)+in_buf[741]*(51)+in_buf[742]*(54)+in_buf[743]*(35)+in_buf[744]*(41)+in_buf[745]*(32)+in_buf[746]*(24)+in_buf[747]*(56)+in_buf[748]*(49)+in_buf[749]*(34)+in_buf[750]*(26)+in_buf[751]*(-2)+in_buf[752]*(2)+in_buf[753]*(5)+in_buf[754]*(1)+in_buf[755]*(4)+in_buf[756]*(3)+in_buf[757]*(3)+in_buf[758]*(-1)+in_buf[759]*(0)+in_buf[760]*(19)+in_buf[761]*(7)+in_buf[762]*(11)+in_buf[763]*(6)+in_buf[764]*(9)+in_buf[765]*(17)+in_buf[766]*(28)+in_buf[767]*(24)+in_buf[768]*(15)+in_buf[769]*(43)+in_buf[770]*(27)+in_buf[771]*(1)+in_buf[772]*(27)+in_buf[773]*(37)+in_buf[774]*(27)+in_buf[775]*(20)+in_buf[776]*(19)+in_buf[777]*(22)+in_buf[778]*(29)+in_buf[779]*(23)+in_buf[780]*(-3)+in_buf[781]*(-2)+in_buf[782]*(-3)+in_buf[783]*(2);
assign in_buf_weight056=in_buf[0]*(-3)+in_buf[1]*(-1)+in_buf[2]*(-1)+in_buf[3]*(1)+in_buf[4]*(0)+in_buf[5]*(-2)+in_buf[6]*(3)+in_buf[7]*(0)+in_buf[8]*(-1)+in_buf[9]*(3)+in_buf[10]*(-1)+in_buf[11]*(2)+in_buf[12]*(16)+in_buf[13]*(8)+in_buf[14]*(-16)+in_buf[15]*(-13)+in_buf[16]*(-3)+in_buf[17]*(0)+in_buf[18]*(3)+in_buf[19]*(2)+in_buf[20]*(0)+in_buf[21]*(1)+in_buf[22]*(3)+in_buf[23]*(-2)+in_buf[24]*(-3)+in_buf[25]*(-3)+in_buf[26]*(-1)+in_buf[27]*(4)+in_buf[28]*(-3)+in_buf[29]*(-1)+in_buf[30]*(0)+in_buf[31]*(-2)+in_buf[32]*(9)+in_buf[33]*(3)+in_buf[34]*(14)+in_buf[35]*(9)+in_buf[36]*(14)+in_buf[37]*(16)+in_buf[38]*(11)+in_buf[39]*(3)+in_buf[40]*(19)+in_buf[41]*(36)+in_buf[42]*(24)+in_buf[43]*(17)+in_buf[44]*(14)+in_buf[45]*(28)+in_buf[46]*(26)+in_buf[47]*(24)+in_buf[48]*(19)+in_buf[49]*(22)+in_buf[50]*(21)+in_buf[51]*(11)+in_buf[52]*(-2)+in_buf[53]*(-3)+in_buf[54]*(3)+in_buf[55]*(3)+in_buf[56]*(2)+in_buf[57]*(-1)+in_buf[58]*(3)+in_buf[59]*(2)+in_buf[60]*(15)+in_buf[61]*(9)+in_buf[62]*(18)+in_buf[63]*(24)+in_buf[64]*(5)+in_buf[65]*(-8)+in_buf[66]*(23)+in_buf[67]*(36)+in_buf[68]*(18)+in_buf[69]*(43)+in_buf[70]*(17)+in_buf[71]*(29)+in_buf[72]*(33)+in_buf[73]*(27)+in_buf[74]*(26)+in_buf[75]*(16)+in_buf[76]*(11)+in_buf[77]*(3)+in_buf[78]*(22)+in_buf[79]*(6)+in_buf[80]*(-3)+in_buf[81]*(-7)+in_buf[82]*(2)+in_buf[83]*(-3)+in_buf[84]*(4)+in_buf[85]*(1)+in_buf[86]*(19)+in_buf[87]*(3)+in_buf[88]*(19)+in_buf[89]*(24)+in_buf[90]*(34)+in_buf[91]*(44)+in_buf[92]*(55)+in_buf[93]*(27)+in_buf[94]*(34)+in_buf[95]*(45)+in_buf[96]*(42)+in_buf[97]*(44)+in_buf[98]*(22)+in_buf[99]*(28)+in_buf[100]*(21)+in_buf[101]*(0)+in_buf[102]*(17)+in_buf[103]*(16)+in_buf[104]*(4)+in_buf[105]*(-6)+in_buf[106]*(-12)+in_buf[107]*(17)+in_buf[108]*(-12)+in_buf[109]*(-38)+in_buf[110]*(-25)+in_buf[111]*(0)+in_buf[112]*(-3)+in_buf[113]*(9)+in_buf[114]*(27)+in_buf[115]*(27)+in_buf[116]*(46)+in_buf[117]*(18)+in_buf[118]*(5)+in_buf[119]*(25)+in_buf[120]*(52)+in_buf[121]*(41)+in_buf[122]*(35)+in_buf[123]*(25)+in_buf[124]*(2)+in_buf[125]*(0)+in_buf[126]*(1)+in_buf[127]*(11)+in_buf[128]*(6)+in_buf[129]*(11)+in_buf[130]*(14)+in_buf[131]*(14)+in_buf[132]*(9)+in_buf[133]*(-2)+in_buf[134]*(8)+in_buf[135]*(-31)+in_buf[136]*(-49)+in_buf[137]*(-12)+in_buf[138]*(12)+in_buf[139]*(17)+in_buf[140]*(0)+in_buf[141]*(1)+in_buf[142]*(15)+in_buf[143]*(39)+in_buf[144]*(39)+in_buf[145]*(0)+in_buf[146]*(-4)+in_buf[147]*(0)+in_buf[148]*(-24)+in_buf[149]*(-17)+in_buf[150]*(-4)+in_buf[151]*(-19)+in_buf[152]*(-15)+in_buf[153]*(-7)+in_buf[154]*(-5)+in_buf[155]*(0)+in_buf[156]*(-7)+in_buf[157]*(0)+in_buf[158]*(3)+in_buf[159]*(25)+in_buf[160]*(32)+in_buf[161]*(23)+in_buf[162]*(11)+in_buf[163]*(-7)+in_buf[164]*(-1)+in_buf[165]*(4)+in_buf[166]*(36)+in_buf[167]*(4)+in_buf[168]*(0)+in_buf[169]*(22)+in_buf[170]*(-2)+in_buf[171]*(20)+in_buf[172]*(16)+in_buf[173]*(-11)+in_buf[174]*(-18)+in_buf[175]*(-22)+in_buf[176]*(-15)+in_buf[177]*(-11)+in_buf[178]*(-7)+in_buf[179]*(-21)+in_buf[180]*(-15)+in_buf[181]*(-5)+in_buf[182]*(-3)+in_buf[183]*(-5)+in_buf[184]*(-7)+in_buf[185]*(-9)+in_buf[186]*(-1)+in_buf[187]*(-8)+in_buf[188]*(-7)+in_buf[189]*(-12)+in_buf[190]*(-9)+in_buf[191]*(1)+in_buf[192]*(2)+in_buf[193]*(16)+in_buf[194]*(44)+in_buf[195]*(32)+in_buf[196]*(1)+in_buf[197]*(20)+in_buf[198]*(-18)+in_buf[199]*(-2)+in_buf[200]*(4)+in_buf[201]*(-2)+in_buf[202]*(-20)+in_buf[203]*(-25)+in_buf[204]*(-13)+in_buf[205]*(-11)+in_buf[206]*(-7)+in_buf[207]*(-5)+in_buf[208]*(0)+in_buf[209]*(-4)+in_buf[210]*(18)+in_buf[211]*(7)+in_buf[212]*(-3)+in_buf[213]*(-6)+in_buf[214]*(0)+in_buf[215]*(2)+in_buf[216]*(-17)+in_buf[217]*(-10)+in_buf[218]*(5)+in_buf[219]*(-9)+in_buf[220]*(-16)+in_buf[221]*(7)+in_buf[222]*(11)+in_buf[223]*(21)+in_buf[224]*(26)+in_buf[225]*(-35)+in_buf[226]*(-11)+in_buf[227]*(13)+in_buf[228]*(-12)+in_buf[229]*(-5)+in_buf[230]*(-6)+in_buf[231]*(-7)+in_buf[232]*(-9)+in_buf[233]*(-5)+in_buf[234]*(-4)+in_buf[235]*(-6)+in_buf[236]*(2)+in_buf[237]*(9)+in_buf[238]*(6)+in_buf[239]*(0)+in_buf[240]*(9)+in_buf[241]*(3)+in_buf[242]*(-2)+in_buf[243]*(0)+in_buf[244]*(-10)+in_buf[245]*(0)+in_buf[246]*(5)+in_buf[247]*(-27)+in_buf[248]*(-38)+in_buf[249]*(3)+in_buf[250]*(5)+in_buf[251]*(19)+in_buf[252]*(-10)+in_buf[253]*(-27)+in_buf[254]*(-27)+in_buf[255]*(4)+in_buf[256]*(-18)+in_buf[257]*(-18)+in_buf[258]*(17)+in_buf[259]*(10)+in_buf[260]*(10)+in_buf[261]*(16)+in_buf[262]*(9)+in_buf[263]*(-2)+in_buf[264]*(-16)+in_buf[265]*(-5)+in_buf[266]*(-4)+in_buf[267]*(1)+in_buf[268]*(9)+in_buf[269]*(-5)+in_buf[270]*(-3)+in_buf[271]*(0)+in_buf[272]*(-7)+in_buf[273]*(-9)+in_buf[274]*(-4)+in_buf[275]*(-2)+in_buf[276]*(-17)+in_buf[277]*(14)+in_buf[278]*(-15)+in_buf[279]*(-25)+in_buf[280]*(-9)+in_buf[281]*(-15)+in_buf[282]*(-10)+in_buf[283]*(26)+in_buf[284]*(-12)+in_buf[285]*(4)+in_buf[286]*(8)+in_buf[287]*(3)+in_buf[288]*(7)+in_buf[289]*(5)+in_buf[290]*(9)+in_buf[291]*(-16)+in_buf[292]*(-22)+in_buf[293]*(-10)+in_buf[294]*(0)+in_buf[295]*(-3)+in_buf[296]*(-1)+in_buf[297]*(8)+in_buf[298]*(4)+in_buf[299]*(-6)+in_buf[300]*(-5)+in_buf[301]*(-18)+in_buf[302]*(-8)+in_buf[303]*(1)+in_buf[304]*(-8)+in_buf[305]*(-28)+in_buf[306]*(-16)+in_buf[307]*(-14)+in_buf[308]*(-10)+in_buf[309]*(-21)+in_buf[310]*(-27)+in_buf[311]*(2)+in_buf[312]*(-14)+in_buf[313]*(-1)+in_buf[314]*(-13)+in_buf[315]*(-16)+in_buf[316]*(-9)+in_buf[317]*(-8)+in_buf[318]*(-12)+in_buf[319]*(-22)+in_buf[320]*(-19)+in_buf[321]*(2)+in_buf[322]*(25)+in_buf[323]*(22)+in_buf[324]*(-3)+in_buf[325]*(0)+in_buf[326]*(5)+in_buf[327]*(1)+in_buf[328]*(-14)+in_buf[329]*(-10)+in_buf[330]*(-22)+in_buf[331]*(-24)+in_buf[332]*(-16)+in_buf[333]*(-13)+in_buf[334]*(18)+in_buf[335]*(-24)+in_buf[336]*(-10)+in_buf[337]*(-19)+in_buf[338]*(-34)+in_buf[339]*(-18)+in_buf[340]*(-9)+in_buf[341]*(2)+in_buf[342]*(-5)+in_buf[343]*(-10)+in_buf[344]*(-26)+in_buf[345]*(-15)+in_buf[346]*(-10)+in_buf[347]*(-14)+in_buf[348]*(9)+in_buf[349]*(20)+in_buf[350]*(29)+in_buf[351]*(3)+in_buf[352]*(-4)+in_buf[353]*(-5)+in_buf[354]*(-11)+in_buf[355]*(-4)+in_buf[356]*(-13)+in_buf[357]*(-2)+in_buf[358]*(-20)+in_buf[359]*(1)+in_buf[360]*(0)+in_buf[361]*(-25)+in_buf[362]*(-26)+in_buf[363]*(-20)+in_buf[364]*(25)+in_buf[365]*(-1)+in_buf[366]*(-27)+in_buf[367]*(-18)+in_buf[368]*(-20)+in_buf[369]*(-18)+in_buf[370]*(-9)+in_buf[371]*(-10)+in_buf[372]*(1)+in_buf[373]*(5)+in_buf[374]*(-1)+in_buf[375]*(0)+in_buf[376]*(17)+in_buf[377]*(24)+in_buf[378]*(5)+in_buf[379]*(-7)+in_buf[380]*(-8)+in_buf[381]*(-5)+in_buf[382]*(6)+in_buf[383]*(4)+in_buf[384]*(-7)+in_buf[385]*(1)+in_buf[386]*(-1)+in_buf[387]*(10)+in_buf[388]*(-16)+in_buf[389]*(12)+in_buf[390]*(4)+in_buf[391]*(17)+in_buf[392]*(13)+in_buf[393]*(-2)+in_buf[394]*(-20)+in_buf[395]*(-5)+in_buf[396]*(-13)+in_buf[397]*(-16)+in_buf[398]*(-1)+in_buf[399]*(0)+in_buf[400]*(9)+in_buf[401]*(1)+in_buf[402]*(-12)+in_buf[403]*(8)+in_buf[404]*(6)+in_buf[405]*(11)+in_buf[406]*(11)+in_buf[407]*(-8)+in_buf[408]*(-6)+in_buf[409]*(4)+in_buf[410]*(5)+in_buf[411]*(-1)+in_buf[412]*(18)+in_buf[413]*(35)+in_buf[414]*(15)+in_buf[415]*(-5)+in_buf[416]*(10)+in_buf[417]*(41)+in_buf[418]*(19)+in_buf[419]*(-8)+in_buf[420]*(10)+in_buf[421]*(12)+in_buf[422]*(15)+in_buf[423]*(-31)+in_buf[424]*(7)+in_buf[425]*(-3)+in_buf[426]*(6)+in_buf[427]*(10)+in_buf[428]*(19)+in_buf[429]*(-2)+in_buf[430]*(-22)+in_buf[431]*(-2)+in_buf[432]*(14)+in_buf[433]*(19)+in_buf[434]*(6)+in_buf[435]*(-16)+in_buf[436]*(0)+in_buf[437]*(2)+in_buf[438]*(-3)+in_buf[439]*(1)+in_buf[440]*(14)+in_buf[441]*(23)+in_buf[442]*(4)+in_buf[443]*(7)+in_buf[444]*(31)+in_buf[445]*(22)+in_buf[446]*(-6)+in_buf[447]*(-1)+in_buf[448]*(0)+in_buf[449]*(19)+in_buf[450]*(25)+in_buf[451]*(13)+in_buf[452]*(17)+in_buf[453]*(22)+in_buf[454]*(8)+in_buf[455]*(1)+in_buf[456]*(4)+in_buf[457]*(0)+in_buf[458]*(-4)+in_buf[459]*(17)+in_buf[460]*(16)+in_buf[461]*(18)+in_buf[462]*(4)+in_buf[463]*(-21)+in_buf[464]*(-14)+in_buf[465]*(-14)+in_buf[466]*(2)+in_buf[467]*(14)+in_buf[468]*(10)+in_buf[469]*(-1)+in_buf[470]*(4)+in_buf[471]*(20)+in_buf[472]*(47)+in_buf[473]*(49)+in_buf[474]*(-4)+in_buf[475]*(-13)+in_buf[476]*(0)+in_buf[477]*(13)+in_buf[478]*(28)+in_buf[479]*(44)+in_buf[480]*(42)+in_buf[481]*(18)+in_buf[482]*(5)+in_buf[483]*(14)+in_buf[484]*(-4)+in_buf[485]*(-13)+in_buf[486]*(10)+in_buf[487]*(5)+in_buf[488]*(7)+in_buf[489]*(18)+in_buf[490]*(-7)+in_buf[491]*(-22)+in_buf[492]*(-2)+in_buf[493]*(8)+in_buf[494]*(2)+in_buf[495]*(22)+in_buf[496]*(-3)+in_buf[497]*(-3)+in_buf[498]*(0)+in_buf[499]*(15)+in_buf[500]*(25)+in_buf[501]*(0)+in_buf[502]*(0)+in_buf[503]*(24)+in_buf[504]*(-35)+in_buf[505]*(17)+in_buf[506]*(25)+in_buf[507]*(51)+in_buf[508]*(28)+in_buf[509]*(10)+in_buf[510]*(11)+in_buf[511]*(-6)+in_buf[512]*(-17)+in_buf[513]*(3)+in_buf[514]*(3)+in_buf[515]*(2)+in_buf[516]*(13)+in_buf[517]*(15)+in_buf[518]*(4)+in_buf[519]*(-7)+in_buf[520]*(7)+in_buf[521]*(8)+in_buf[522]*(4)+in_buf[523]*(12)+in_buf[524]*(10)+in_buf[525]*(7)+in_buf[526]*(0)+in_buf[527]*(27)+in_buf[528]*(34)+in_buf[529]*(22)+in_buf[530]*(-26)+in_buf[531]*(-9)+in_buf[532]*(20)+in_buf[533]*(-38)+in_buf[534]*(-15)+in_buf[535]*(42)+in_buf[536]*(5)+in_buf[537]*(19)+in_buf[538]*(6)+in_buf[539]*(5)+in_buf[540]*(-2)+in_buf[541]*(19)+in_buf[542]*(26)+in_buf[543]*(25)+in_buf[544]*(26)+in_buf[545]*(25)+in_buf[546]*(14)+in_buf[547]*(14)+in_buf[548]*(19)+in_buf[549]*(13)+in_buf[550]*(28)+in_buf[551]*(17)+in_buf[552]*(16)+in_buf[553]*(24)+in_buf[554]*(21)+in_buf[555]*(47)+in_buf[556]*(53)+in_buf[557]*(37)+in_buf[558]*(-5)+in_buf[559]*(-8)+in_buf[560]*(0)+in_buf[561]*(-2)+in_buf[562]*(-15)+in_buf[563]*(20)+in_buf[564]*(10)+in_buf[565]*(-14)+in_buf[566]*(-2)+in_buf[567]*(12)+in_buf[568]*(6)+in_buf[569]*(31)+in_buf[570]*(26)+in_buf[571]*(31)+in_buf[572]*(24)+in_buf[573]*(23)+in_buf[574]*(30)+in_buf[575]*(20)+in_buf[576]*(12)+in_buf[577]*(9)+in_buf[578]*(30)+in_buf[579]*(17)+in_buf[580]*(36)+in_buf[581]*(35)+in_buf[582]*(28)+in_buf[583]*(23)+in_buf[584]*(28)+in_buf[585]*(21)+in_buf[586]*(15)+in_buf[587]*(10)+in_buf[588]*(10)+in_buf[589]*(8)+in_buf[590]*(0)+in_buf[591]*(24)+in_buf[592]*(-10)+in_buf[593]*(-44)+in_buf[594]*(-6)+in_buf[595]*(9)+in_buf[596]*(15)+in_buf[597]*(3)+in_buf[598]*(1)+in_buf[599]*(17)+in_buf[600]*(14)+in_buf[601]*(22)+in_buf[602]*(23)+in_buf[603]*(14)+in_buf[604]*(0)+in_buf[605]*(3)+in_buf[606]*(11)+in_buf[607]*(15)+in_buf[608]*(29)+in_buf[609]*(-1)+in_buf[610]*(27)+in_buf[611]*(4)+in_buf[612]*(-14)+in_buf[613]*(3)+in_buf[614]*(-4)+in_buf[615]*(-5)+in_buf[616]*(11)+in_buf[617]*(28)+in_buf[618]*(11)+in_buf[619]*(15)+in_buf[620]*(0)+in_buf[621]*(-12)+in_buf[622]*(-19)+in_buf[623]*(-9)+in_buf[624]*(-10)+in_buf[625]*(-2)+in_buf[626]*(-7)+in_buf[627]*(9)+in_buf[628]*(-3)+in_buf[629]*(13)+in_buf[630]*(7)+in_buf[631]*(5)+in_buf[632]*(1)+in_buf[633]*(8)+in_buf[634]*(10)+in_buf[635]*(13)+in_buf[636]*(16)+in_buf[637]*(6)+in_buf[638]*(33)+in_buf[639]*(8)+in_buf[640]*(-16)+in_buf[641]*(20)+in_buf[642]*(18)+in_buf[643]*(-1)+in_buf[644]*(2)+in_buf[645]*(2)+in_buf[646]*(39)+in_buf[647]*(42)+in_buf[648]*(1)+in_buf[649]*(12)+in_buf[650]*(3)+in_buf[651]*(-5)+in_buf[652]*(2)+in_buf[653]*(12)+in_buf[654]*(6)+in_buf[655]*(20)+in_buf[656]*(8)+in_buf[657]*(10)+in_buf[658]*(2)+in_buf[659]*(8)+in_buf[660]*(3)+in_buf[661]*(11)+in_buf[662]*(15)+in_buf[663]*(-6)+in_buf[664]*(2)+in_buf[665]*(7)+in_buf[666]*(16)+in_buf[667]*(8)+in_buf[668]*(-8)+in_buf[669]*(12)+in_buf[670]*(23)+in_buf[671]*(0)+in_buf[672]*(1)+in_buf[673]*(0)+in_buf[674]*(11)+in_buf[675]*(26)+in_buf[676]*(7)+in_buf[677]*(-7)+in_buf[678]*(8)+in_buf[679]*(9)+in_buf[680]*(8)+in_buf[681]*(11)+in_buf[682]*(9)+in_buf[683]*(0)+in_buf[684]*(10)+in_buf[685]*(-6)+in_buf[686]*(5)+in_buf[687]*(-9)+in_buf[688]*(1)+in_buf[689]*(-2)+in_buf[690]*(-6)+in_buf[691]*(-32)+in_buf[692]*(-6)+in_buf[693]*(-11)+in_buf[694]*(1)+in_buf[695]*(28)+in_buf[696]*(6)+in_buf[697]*(-6)+in_buf[698]*(-3)+in_buf[699]*(0)+in_buf[700]*(2)+in_buf[701]*(1)+in_buf[702]*(19)+in_buf[703]*(-17)+in_buf[704]*(-13)+in_buf[705]*(-3)+in_buf[706]*(8)+in_buf[707]*(6)+in_buf[708]*(0)+in_buf[709]*(4)+in_buf[710]*(11)+in_buf[711]*(5)+in_buf[712]*(0)+in_buf[713]*(10)+in_buf[714]*(-11)+in_buf[715]*(-8)+in_buf[716]*(0)+in_buf[717]*(-21)+in_buf[718]*(-21)+in_buf[719]*(10)+in_buf[720]*(5)+in_buf[721]*(-15)+in_buf[722]*(-17)+in_buf[723]*(13)+in_buf[724]*(9)+in_buf[725]*(-1)+in_buf[726]*(2)+in_buf[727]*(-3)+in_buf[728]*(4)+in_buf[729]*(2)+in_buf[730]*(0)+in_buf[731]*(-7)+in_buf[732]*(26)+in_buf[733]*(31)+in_buf[734]*(-1)+in_buf[735]*(-27)+in_buf[736]*(-32)+in_buf[737]*(-31)+in_buf[738]*(-3)+in_buf[739]*(8)+in_buf[740]*(16)+in_buf[741]*(8)+in_buf[742]*(-8)+in_buf[743]*(-12)+in_buf[744]*(22)+in_buf[745]*(22)+in_buf[746]*(17)+in_buf[747]*(-4)+in_buf[748]*(4)+in_buf[749]*(2)+in_buf[750]*(7)+in_buf[751]*(8)+in_buf[752]*(23)+in_buf[753]*(1)+in_buf[754]*(2)+in_buf[755]*(-2)+in_buf[756]*(3)+in_buf[757]*(2)+in_buf[758]*(2)+in_buf[759]*(3)+in_buf[760]*(-14)+in_buf[761]*(-18)+in_buf[762]*(16)+in_buf[763]*(17)+in_buf[764]*(11)+in_buf[765]*(-10)+in_buf[766]*(-26)+in_buf[767]*(-5)+in_buf[768]*(10)+in_buf[769]*(-22)+in_buf[770]*(-1)+in_buf[771]*(14)+in_buf[772]*(0)+in_buf[773]*(-21)+in_buf[774]*(-11)+in_buf[775]*(6)+in_buf[776]*(0)+in_buf[777]*(-15)+in_buf[778]*(-12)+in_buf[779]*(-19)+in_buf[780]*(1)+in_buf[781]*(0)+in_buf[782]*(1)+in_buf[783]*(2);
assign in_buf_weight057=in_buf[0]*(0)+in_buf[1]*(3)+in_buf[2]*(4)+in_buf[3]*(-3)+in_buf[4]*(-2)+in_buf[5]*(0)+in_buf[6]*(4)+in_buf[7]*(-2)+in_buf[8]*(-2)+in_buf[9]*(1)+in_buf[10]*(-1)+in_buf[11]*(1)+in_buf[12]*(8)+in_buf[13]*(7)+in_buf[14]*(-4)+in_buf[15]*(-3)+in_buf[16]*(4)+in_buf[17]*(4)+in_buf[18]*(3)+in_buf[19]*(1)+in_buf[20]*(1)+in_buf[21]*(-2)+in_buf[22]*(-3)+in_buf[23]*(0)+in_buf[24]*(-3)+in_buf[25]*(-1)+in_buf[26]*(3)+in_buf[27]*(0)+in_buf[28]*(0)+in_buf[29]*(-1)+in_buf[30]*(2)+in_buf[31]*(4)+in_buf[32]*(5)+in_buf[33]*(4)+in_buf[34]*(14)+in_buf[35]*(11)+in_buf[36]*(15)+in_buf[37]*(8)+in_buf[38]*(17)+in_buf[39]*(33)+in_buf[40]*(42)+in_buf[41]*(31)+in_buf[42]*(-6)+in_buf[43]*(27)+in_buf[44]*(14)+in_buf[45]*(28)+in_buf[46]*(14)+in_buf[47]*(9)+in_buf[48]*(16)+in_buf[49]*(13)+in_buf[50]*(6)+in_buf[51]*(10)+in_buf[52]*(-1)+in_buf[53]*(3)+in_buf[54]*(3)+in_buf[55]*(4)+in_buf[56]*(2)+in_buf[57]*(-3)+in_buf[58]*(17)+in_buf[59]*(26)+in_buf[60]*(30)+in_buf[61]*(11)+in_buf[62]*(16)+in_buf[63]*(28)+in_buf[64]*(16)+in_buf[65]*(3)+in_buf[66]*(21)+in_buf[67]*(60)+in_buf[68]*(32)+in_buf[69]*(-5)+in_buf[70]*(-12)+in_buf[71]*(0)+in_buf[72]*(7)+in_buf[73]*(5)+in_buf[74]*(0)+in_buf[75]*(2)+in_buf[76]*(0)+in_buf[77]*(-3)+in_buf[78]*(8)+in_buf[79]*(-4)+in_buf[80]*(-3)+in_buf[81]*(0)+in_buf[82]*(0)+in_buf[83]*(1)+in_buf[84]*(4)+in_buf[85]*(-3)+in_buf[86]*(12)+in_buf[87]*(37)+in_buf[88]*(31)+in_buf[89]*(2)+in_buf[90]*(28)+in_buf[91]*(24)+in_buf[92]*(36)+in_buf[93]*(52)+in_buf[94]*(37)+in_buf[95]*(19)+in_buf[96]*(24)+in_buf[97]*(44)+in_buf[98]*(38)+in_buf[99]*(18)+in_buf[100]*(5)+in_buf[101]*(0)+in_buf[102]*(2)+in_buf[103]*(12)+in_buf[104]*(-10)+in_buf[105]*(-4)+in_buf[106]*(0)+in_buf[107]*(8)+in_buf[108]*(-1)+in_buf[109]*(9)+in_buf[110]*(3)+in_buf[111]*(0)+in_buf[112]*(4)+in_buf[113]*(1)+in_buf[114]*(1)+in_buf[115]*(0)+in_buf[116]*(39)+in_buf[117]*(11)+in_buf[118]*(13)+in_buf[119]*(5)+in_buf[120]*(15)+in_buf[121]*(33)+in_buf[122]*(18)+in_buf[123]*(4)+in_buf[124]*(13)+in_buf[125]*(27)+in_buf[126]*(28)+in_buf[127]*(22)+in_buf[128]*(21)+in_buf[129]*(14)+in_buf[130]*(14)+in_buf[131]*(9)+in_buf[132]*(26)+in_buf[133]*(5)+in_buf[134]*(-5)+in_buf[135]*(-22)+in_buf[136]*(-45)+in_buf[137]*(-30)+in_buf[138]*(-8)+in_buf[139]*(-1)+in_buf[140]*(0)+in_buf[141]*(-1)+in_buf[142]*(0)+in_buf[143]*(-38)+in_buf[144]*(-18)+in_buf[145]*(-17)+in_buf[146]*(3)+in_buf[147]*(-1)+in_buf[148]*(22)+in_buf[149]*(10)+in_buf[150]*(0)+in_buf[151]*(-14)+in_buf[152]*(-9)+in_buf[153]*(1)+in_buf[154]*(2)+in_buf[155]*(-7)+in_buf[156]*(-3)+in_buf[157]*(0)+in_buf[158]*(1)+in_buf[159]*(0)+in_buf[160]*(-10)+in_buf[161]*(-14)+in_buf[162]*(-12)+in_buf[163]*(-33)+in_buf[164]*(-45)+in_buf[165]*(-46)+in_buf[166]*(-4)+in_buf[167]*(1)+in_buf[168]*(0)+in_buf[169]*(-2)+in_buf[170]*(15)+in_buf[171]*(-3)+in_buf[172]*(21)+in_buf[173]*(27)+in_buf[174]*(-9)+in_buf[175]*(-11)+in_buf[176]*(1)+in_buf[177]*(-25)+in_buf[178]*(-24)+in_buf[179]*(8)+in_buf[180]*(8)+in_buf[181]*(3)+in_buf[182]*(0)+in_buf[183]*(-7)+in_buf[184]*(-29)+in_buf[185]*(-21)+in_buf[186]*(-6)+in_buf[187]*(-14)+in_buf[188]*(-13)+in_buf[189]*(11)+in_buf[190]*(-13)+in_buf[191]*(-28)+in_buf[192]*(-19)+in_buf[193]*(-41)+in_buf[194]*(-33)+in_buf[195]*(-13)+in_buf[196]*(6)+in_buf[197]*(27)+in_buf[198]*(0)+in_buf[199]*(2)+in_buf[200]*(11)+in_buf[201]*(17)+in_buf[202]*(-2)+in_buf[203]*(16)+in_buf[204]*(-3)+in_buf[205]*(0)+in_buf[206]*(12)+in_buf[207]*(22)+in_buf[208]*(12)+in_buf[209]*(0)+in_buf[210]*(-1)+in_buf[211]*(-8)+in_buf[212]*(-10)+in_buf[213]*(-10)+in_buf[214]*(1)+in_buf[215]*(-2)+in_buf[216]*(-5)+in_buf[217]*(-6)+in_buf[218]*(-7)+in_buf[219]*(-22)+in_buf[220]*(-2)+in_buf[221]*(-34)+in_buf[222]*(-30)+in_buf[223]*(0)+in_buf[224]*(8)+in_buf[225]*(40)+in_buf[226]*(6)+in_buf[227]*(1)+in_buf[228]*(16)+in_buf[229]*(14)+in_buf[230]*(14)+in_buf[231]*(11)+in_buf[232]*(13)+in_buf[233]*(11)+in_buf[234]*(14)+in_buf[235]*(16)+in_buf[236]*(21)+in_buf[237]*(-2)+in_buf[238]*(-15)+in_buf[239]*(-13)+in_buf[240]*(-17)+in_buf[241]*(-10)+in_buf[242]*(-7)+in_buf[243]*(-12)+in_buf[244]*(-1)+in_buf[245]*(-9)+in_buf[246]*(2)+in_buf[247]*(9)+in_buf[248]*(-6)+in_buf[249]*(-24)+in_buf[250]*(-46)+in_buf[251]*(-14)+in_buf[252]*(22)+in_buf[253]*(38)+in_buf[254]*(0)+in_buf[255]*(16)+in_buf[256]*(49)+in_buf[257]*(30)+in_buf[258]*(13)+in_buf[259]*(22)+in_buf[260]*(10)+in_buf[261]*(7)+in_buf[262]*(21)+in_buf[263]*(31)+in_buf[264]*(23)+in_buf[265]*(-2)+in_buf[266]*(-19)+in_buf[267]*(-22)+in_buf[268]*(-13)+in_buf[269]*(-7)+in_buf[270]*(1)+in_buf[271]*(-9)+in_buf[272]*(2)+in_buf[273]*(12)+in_buf[274]*(18)+in_buf[275]*(26)+in_buf[276]*(16)+in_buf[277]*(0)+in_buf[278]*(-32)+in_buf[279]*(-2)+in_buf[280]*(21)+in_buf[281]*(31)+in_buf[282]*(40)+in_buf[283]*(0)+in_buf[284]*(39)+in_buf[285]*(22)+in_buf[286]*(6)+in_buf[287]*(0)+in_buf[288]*(7)+in_buf[289]*(25)+in_buf[290]*(40)+in_buf[291]*(43)+in_buf[292]*(17)+in_buf[293]*(-7)+in_buf[294]*(-20)+in_buf[295]*(-13)+in_buf[296]*(5)+in_buf[297]*(17)+in_buf[298]*(13)+in_buf[299]*(16)+in_buf[300]*(17)+in_buf[301]*(26)+in_buf[302]*(28)+in_buf[303]*(21)+in_buf[304]*(49)+in_buf[305]*(13)+in_buf[306]*(0)+in_buf[307]*(-10)+in_buf[308]*(19)+in_buf[309]*(50)+in_buf[310]*(37)+in_buf[311]*(16)+in_buf[312]*(17)+in_buf[313]*(-2)+in_buf[314]*(4)+in_buf[315]*(-4)+in_buf[316]*(1)+in_buf[317]*(31)+in_buf[318]*(42)+in_buf[319]*(45)+in_buf[320]*(12)+in_buf[321]*(-20)+in_buf[322]*(-33)+in_buf[323]*(-17)+in_buf[324]*(11)+in_buf[325]*(22)+in_buf[326]*(33)+in_buf[327]*(18)+in_buf[328]*(13)+in_buf[329]*(15)+in_buf[330]*(19)+in_buf[331]*(31)+in_buf[332]*(55)+in_buf[333]*(3)+in_buf[334]*(0)+in_buf[335]*(0)+in_buf[336]*(26)+in_buf[337]*(27)+in_buf[338]*(5)+in_buf[339]*(21)+in_buf[340]*(3)+in_buf[341]*(-2)+in_buf[342]*(4)+in_buf[343]*(15)+in_buf[344]*(22)+in_buf[345]*(43)+in_buf[346]*(48)+in_buf[347]*(32)+in_buf[348]*(-11)+in_buf[349]*(-33)+in_buf[350]*(-21)+in_buf[351]*(-5)+in_buf[352]*(19)+in_buf[353]*(14)+in_buf[354]*(22)+in_buf[355]*(1)+in_buf[356]*(21)+in_buf[357]*(11)+in_buf[358]*(28)+in_buf[359]*(36)+in_buf[360]*(42)+in_buf[361]*(-11)+in_buf[362]*(7)+in_buf[363]*(0)+in_buf[364]*(1)+in_buf[365]*(12)+in_buf[366]*(33)+in_buf[367]*(31)+in_buf[368]*(7)+in_buf[369]*(13)+in_buf[370]*(19)+in_buf[371]*(8)+in_buf[372]*(21)+in_buf[373]*(39)+in_buf[374]*(24)+in_buf[375]*(2)+in_buf[376]*(-36)+in_buf[377]*(-34)+in_buf[378]*(-10)+in_buf[379]*(-12)+in_buf[380]*(-5)+in_buf[381]*(-5)+in_buf[382]*(2)+in_buf[383]*(0)+in_buf[384]*(4)+in_buf[385]*(15)+in_buf[386]*(9)+in_buf[387]*(32)+in_buf[388]*(30)+in_buf[389]*(0)+in_buf[390]*(-21)+in_buf[391]*(-13)+in_buf[392]*(6)+in_buf[393]*(12)+in_buf[394]*(36)+in_buf[395]*(13)+in_buf[396]*(-13)+in_buf[397]*(22)+in_buf[398]*(4)+in_buf[399]*(5)+in_buf[400]*(25)+in_buf[401]*(34)+in_buf[402]*(28)+in_buf[403]*(-6)+in_buf[404]*(-37)+in_buf[405]*(-32)+in_buf[406]*(-15)+in_buf[407]*(-8)+in_buf[408]*(-15)+in_buf[409]*(-17)+in_buf[410]*(-7)+in_buf[411]*(-10)+in_buf[412]*(-8)+in_buf[413]*(-3)+in_buf[414]*(15)+in_buf[415]*(58)+in_buf[416]*(58)+in_buf[417]*(-1)+in_buf[418]*(-17)+in_buf[419]*(-6)+in_buf[420]*(8)+in_buf[421]*(-1)+in_buf[422]*(22)+in_buf[423]*(21)+in_buf[424]*(-21)+in_buf[425]*(13)+in_buf[426]*(15)+in_buf[427]*(24)+in_buf[428]*(19)+in_buf[429]*(12)+in_buf[430]*(8)+in_buf[431]*(-15)+in_buf[432]*(-26)+in_buf[433]*(-30)+in_buf[434]*(-16)+in_buf[435]*(-6)+in_buf[436]*(-24)+in_buf[437]*(-13)+in_buf[438]*(-16)+in_buf[439]*(-17)+in_buf[440]*(-7)+in_buf[441]*(6)+in_buf[442]*(22)+in_buf[443]*(38)+in_buf[444]*(21)+in_buf[445]*(11)+in_buf[446]*(-35)+in_buf[447]*(-33)+in_buf[448]*(7)+in_buf[449]*(0)+in_buf[450]*(14)+in_buf[451]*(25)+in_buf[452]*(7)+in_buf[453]*(19)+in_buf[454]*(7)+in_buf[455]*(22)+in_buf[456]*(39)+in_buf[457]*(27)+in_buf[458]*(3)+in_buf[459]*(-17)+in_buf[460]*(-35)+in_buf[461]*(-44)+in_buf[462]*(-14)+in_buf[463]*(-13)+in_buf[464]*(-35)+in_buf[465]*(-32)+in_buf[466]*(-36)+in_buf[467]*(-12)+in_buf[468]*(-12)+in_buf[469]*(5)+in_buf[470]*(21)+in_buf[471]*(26)+in_buf[472]*(23)+in_buf[473]*(9)+in_buf[474]*(-43)+in_buf[475]*(-30)+in_buf[476]*(-3)+in_buf[477]*(-3)+in_buf[478]*(18)+in_buf[479]*(15)+in_buf[480]*(21)+in_buf[481]*(28)+in_buf[482]*(2)+in_buf[483]*(11)+in_buf[484]*(12)+in_buf[485]*(2)+in_buf[486]*(-7)+in_buf[487]*(-2)+in_buf[488]*(-25)+in_buf[489]*(-27)+in_buf[490]*(0)+in_buf[491]*(-26)+in_buf[492]*(-38)+in_buf[493]*(-29)+in_buf[494]*(-14)+in_buf[495]*(-10)+in_buf[496]*(0)+in_buf[497]*(17)+in_buf[498]*(35)+in_buf[499]*(42)+in_buf[500]*(5)+in_buf[501]*(5)+in_buf[502]*(-31)+in_buf[503]*(-14)+in_buf[504]*(9)+in_buf[505]*(-1)+in_buf[506]*(17)+in_buf[507]*(6)+in_buf[508]*(4)+in_buf[509]*(15)+in_buf[510]*(-3)+in_buf[511]*(0)+in_buf[512]*(-1)+in_buf[513]*(-1)+in_buf[514]*(2)+in_buf[515]*(-1)+in_buf[516]*(-10)+in_buf[517]*(-22)+in_buf[518]*(-12)+in_buf[519]*(-16)+in_buf[520]*(-11)+in_buf[521]*(-19)+in_buf[522]*(0)+in_buf[523]*(-1)+in_buf[524]*(16)+in_buf[525]*(31)+in_buf[526]*(25)+in_buf[527]*(19)+in_buf[528]*(1)+in_buf[529]*(5)+in_buf[530]*(-33)+in_buf[531]*(-29)+in_buf[532]*(3)+in_buf[533]*(40)+in_buf[534]*(26)+in_buf[535]*(18)+in_buf[536]*(16)+in_buf[537]*(9)+in_buf[538]*(8)+in_buf[539]*(4)+in_buf[540]*(-4)+in_buf[541]*(5)+in_buf[542]*(2)+in_buf[543]*(16)+in_buf[544]*(0)+in_buf[545]*(-24)+in_buf[546]*(-17)+in_buf[547]*(-15)+in_buf[548]*(-17)+in_buf[549]*(-12)+in_buf[550]*(0)+in_buf[551]*(13)+in_buf[552]*(34)+in_buf[553]*(25)+in_buf[554]*(17)+in_buf[555]*(2)+in_buf[556]*(3)+in_buf[557]*(-23)+in_buf[558]*(-39)+in_buf[559]*(-22)+in_buf[560]*(2)+in_buf[561]*(7)+in_buf[562]*(7)+in_buf[563]*(13)+in_buf[564]*(21)+in_buf[565]*(-11)+in_buf[566]*(-1)+in_buf[567]*(9)+in_buf[568]*(5)+in_buf[569]*(13)+in_buf[570]*(11)+in_buf[571]*(15)+in_buf[572]*(18)+in_buf[573]*(-15)+in_buf[574]*(-6)+in_buf[575]*(-11)+in_buf[576]*(-15)+in_buf[577]*(-2)+in_buf[578]*(13)+in_buf[579]*(22)+in_buf[580]*(12)+in_buf[581]*(4)+in_buf[582]*(17)+in_buf[583]*(-8)+in_buf[584]*(-9)+in_buf[585]*(-40)+in_buf[586]*(-24)+in_buf[587]*(-5)+in_buf[588]*(0)+in_buf[589]*(-3)+in_buf[590]*(-12)+in_buf[591]*(-14)+in_buf[592]*(16)+in_buf[593]*(-23)+in_buf[594]*(-13)+in_buf[595]*(-17)+in_buf[596]*(-2)+in_buf[597]*(6)+in_buf[598]*(13)+in_buf[599]*(22)+in_buf[600]*(12)+in_buf[601]*(6)+in_buf[602]*(2)+in_buf[603]*(0)+in_buf[604]*(1)+in_buf[605]*(12)+in_buf[606]*(23)+in_buf[607]*(31)+in_buf[608]*(21)+in_buf[609]*(14)+in_buf[610]*(14)+in_buf[611]*(-14)+in_buf[612]*(-32)+in_buf[613]*(-17)+in_buf[614]*(22)+in_buf[615]*(3)+in_buf[616]*(0)+in_buf[617]*(0)+in_buf[618]*(-6)+in_buf[619]*(-15)+in_buf[620]*(-11)+in_buf[621]*(-13)+in_buf[622]*(-35)+in_buf[623]*(-28)+in_buf[624]*(-6)+in_buf[625]*(-8)+in_buf[626]*(-18)+in_buf[627]*(-16)+in_buf[628]*(-2)+in_buf[629]*(13)+in_buf[630]*(11)+in_buf[631]*(22)+in_buf[632]*(20)+in_buf[633]*(26)+in_buf[634]*(22)+in_buf[635]*(38)+in_buf[636]*(7)+in_buf[637]*(6)+in_buf[638]*(3)+in_buf[639]*(-17)+in_buf[640]*(-61)+in_buf[641]*(-33)+in_buf[642]*(40)+in_buf[643]*(6)+in_buf[644]*(2)+in_buf[645]*(-1)+in_buf[646]*(-1)+in_buf[647]*(-4)+in_buf[648]*(-28)+in_buf[649]*(-2)+in_buf[650]*(0)+in_buf[651]*(-16)+in_buf[652]*(-10)+in_buf[653]*(-2)+in_buf[654]*(-14)+in_buf[655]*(-17)+in_buf[656]*(-5)+in_buf[657]*(0)+in_buf[658]*(18)+in_buf[659]*(11)+in_buf[660]*(9)+in_buf[661]*(16)+in_buf[662]*(7)+in_buf[663]*(9)+in_buf[664]*(-22)+in_buf[665]*(-7)+in_buf[666]*(-16)+in_buf[667]*(-43)+in_buf[668]*(-50)+in_buf[669]*(-18)+in_buf[670]*(6)+in_buf[671]*(4)+in_buf[672]*(0)+in_buf[673]*(-1)+in_buf[674]*(-2)+in_buf[675]*(0)+in_buf[676]*(14)+in_buf[677]*(2)+in_buf[678]*(4)+in_buf[679]*(24)+in_buf[680]*(1)+in_buf[681]*(5)+in_buf[682]*(-2)+in_buf[683]*(-9)+in_buf[684]*(-8)+in_buf[685]*(8)+in_buf[686]*(9)+in_buf[687]*(6)+in_buf[688]*(-9)+in_buf[689]*(15)+in_buf[690]*(8)+in_buf[691]*(-3)+in_buf[692]*(-20)+in_buf[693]*(-1)+in_buf[694]*(8)+in_buf[695]*(-38)+in_buf[696]*(-31)+in_buf[697]*(-13)+in_buf[698]*(1)+in_buf[699]*(0)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(-26)+in_buf[703]*(9)+in_buf[704]*(5)+in_buf[705]*(-15)+in_buf[706]*(-1)+in_buf[707]*(0)+in_buf[708]*(0)+in_buf[709]*(-1)+in_buf[710]*(-13)+in_buf[711]*(6)+in_buf[712]*(1)+in_buf[713]*(4)+in_buf[714]*(6)+in_buf[715]*(10)+in_buf[716]*(18)+in_buf[717]*(25)+in_buf[718]*(13)+in_buf[719]*(5)+in_buf[720]*(11)+in_buf[721]*(31)+in_buf[722]*(27)+in_buf[723]*(1)+in_buf[724]*(9)+in_buf[725]*(4)+in_buf[726]*(-3)+in_buf[727]*(1)+in_buf[728]*(3)+in_buf[729]*(4)+in_buf[730]*(0)+in_buf[731]*(-3)+in_buf[732]*(-6)+in_buf[733]*(-10)+in_buf[734]*(-3)+in_buf[735]*(0)+in_buf[736]*(-5)+in_buf[737]*(11)+in_buf[738]*(-2)+in_buf[739]*(5)+in_buf[740]*(-7)+in_buf[741]*(-10)+in_buf[742]*(-6)+in_buf[743]*(0)+in_buf[744]*(4)+in_buf[745]*(2)+in_buf[746]*(6)+in_buf[747]*(28)+in_buf[748]*(6)+in_buf[749]*(0)+in_buf[750]*(3)+in_buf[751]*(-11)+in_buf[752]*(-30)+in_buf[753]*(12)+in_buf[754]*(-1)+in_buf[755]*(2)+in_buf[756]*(0)+in_buf[757]*(0)+in_buf[758]*(0)+in_buf[759]*(0)+in_buf[760]*(28)+in_buf[761]*(31)+in_buf[762]*(17)+in_buf[763]*(7)+in_buf[764]*(18)+in_buf[765]*(31)+in_buf[766]*(19)+in_buf[767]*(28)+in_buf[768]*(17)+in_buf[769]*(40)+in_buf[770]*(4)+in_buf[771]*(-11)+in_buf[772]*(16)+in_buf[773]*(31)+in_buf[774]*(7)+in_buf[775]*(-19)+in_buf[776]*(2)+in_buf[777]*(24)+in_buf[778]*(22)+in_buf[779]*(33)+in_buf[780]*(-2)+in_buf[781]*(4)+in_buf[782]*(-1)+in_buf[783]*(-2);
assign in_buf_weight058=in_buf[0]*(4)+in_buf[1]*(-3)+in_buf[2]*(-1)+in_buf[3]*(4)+in_buf[4]*(2)+in_buf[5]*(-2)+in_buf[6]*(-1)+in_buf[7]*(2)+in_buf[8]*(-2)+in_buf[9]*(2)+in_buf[10]*(-1)+in_buf[11]*(1)+in_buf[12]*(10)+in_buf[13]*(10)+in_buf[14]*(-21)+in_buf[15]*(-11)+in_buf[16]*(4)+in_buf[17]*(2)+in_buf[18]*(3)+in_buf[19]*(0)+in_buf[20]*(1)+in_buf[21]*(3)+in_buf[22]*(1)+in_buf[23]*(-2)+in_buf[24]*(-3)+in_buf[25]*(-2)+in_buf[26]*(-1)+in_buf[27]*(4)+in_buf[28]*(-1)+in_buf[29]*(0)+in_buf[30]*(2)+in_buf[31]*(3)+in_buf[32]*(1)+in_buf[33]*(6)+in_buf[34]*(4)+in_buf[35]*(14)+in_buf[36]*(17)+in_buf[37]*(5)+in_buf[38]*(-7)+in_buf[39]*(12)+in_buf[40]*(22)+in_buf[41]*(32)+in_buf[42]*(-16)+in_buf[43]*(1)+in_buf[44]*(21)+in_buf[45]*(34)+in_buf[46]*(27)+in_buf[47]*(32)+in_buf[48]*(48)+in_buf[49]*(33)+in_buf[50]*(21)+in_buf[51]*(7)+in_buf[52]*(0)+in_buf[53]*(-1)+in_buf[54]*(-2)+in_buf[55]*(2)+in_buf[56]*(4)+in_buf[57]*(2)+in_buf[58]*(12)+in_buf[59]*(10)+in_buf[60]*(19)+in_buf[61]*(1)+in_buf[62]*(11)+in_buf[63]*(21)+in_buf[64]*(21)+in_buf[65]*(-3)+in_buf[66]*(-28)+in_buf[67]*(7)+in_buf[68]*(14)+in_buf[69]*(-21)+in_buf[70]*(3)+in_buf[71]*(-14)+in_buf[72]*(-22)+in_buf[73]*(-9)+in_buf[74]*(1)+in_buf[75]*(32)+in_buf[76]*(26)+in_buf[77]*(34)+in_buf[78]*(31)+in_buf[79]*(-2)+in_buf[80]*(-3)+in_buf[81]*(-1)+in_buf[82]*(4)+in_buf[83]*(-1)+in_buf[84]*(3)+in_buf[85]*(3)+in_buf[86]*(-22)+in_buf[87]*(19)+in_buf[88]*(2)+in_buf[89]*(28)+in_buf[90]*(22)+in_buf[91]*(44)+in_buf[92]*(42)+in_buf[93]*(2)+in_buf[94]*(10)+in_buf[95]*(45)+in_buf[96]*(24)+in_buf[97]*(28)+in_buf[98]*(43)+in_buf[99]*(13)+in_buf[100]*(1)+in_buf[101]*(-3)+in_buf[102]*(-13)+in_buf[103]*(-6)+in_buf[104]*(11)+in_buf[105]*(13)+in_buf[106]*(-1)+in_buf[107]*(9)+in_buf[108]*(8)+in_buf[109]*(-9)+in_buf[110]*(-16)+in_buf[111]*(5)+in_buf[112]*(3)+in_buf[113]*(3)+in_buf[114]*(5)+in_buf[115]*(30)+in_buf[116]*(37)+in_buf[117]*(22)+in_buf[118]*(7)+in_buf[119]*(16)+in_buf[120]*(32)+in_buf[121]*(14)+in_buf[122]*(20)+in_buf[123]*(20)+in_buf[124]*(7)+in_buf[125]*(-2)+in_buf[126]*(-3)+in_buf[127]*(-13)+in_buf[128]*(-7)+in_buf[129]*(-8)+in_buf[130]*(-10)+in_buf[131]*(1)+in_buf[132]*(0)+in_buf[133]*(-13)+in_buf[134]*(-17)+in_buf[135]*(-50)+in_buf[136]*(-32)+in_buf[137]*(-25)+in_buf[138]*(-3)+in_buf[139]*(28)+in_buf[140]*(4)+in_buf[141]*(-2)+in_buf[142]*(21)+in_buf[143]*(17)+in_buf[144]*(18)+in_buf[145]*(16)+in_buf[146]*(19)+in_buf[147]*(23)+in_buf[148]*(13)+in_buf[149]*(18)+in_buf[150]*(12)+in_buf[151]*(-4)+in_buf[152]*(7)+in_buf[153]*(4)+in_buf[154]*(5)+in_buf[155]*(-2)+in_buf[156]*(-6)+in_buf[157]*(-6)+in_buf[158]*(-3)+in_buf[159]*(0)+in_buf[160]*(-32)+in_buf[161]*(-44)+in_buf[162]*(-41)+in_buf[163]*(-29)+in_buf[164]*(-11)+in_buf[165]*(17)+in_buf[166]*(9)+in_buf[167]*(12)+in_buf[168]*(0)+in_buf[169]*(24)+in_buf[170]*(12)+in_buf[171]*(21)+in_buf[172]*(29)+in_buf[173]*(27)+in_buf[174]*(22)+in_buf[175]*(10)+in_buf[176]*(18)+in_buf[177]*(15)+in_buf[178]*(10)+in_buf[179]*(-5)+in_buf[180]*(-3)+in_buf[181]*(9)+in_buf[182]*(0)+in_buf[183]*(3)+in_buf[184]*(7)+in_buf[185]*(0)+in_buf[186]*(-10)+in_buf[187]*(-8)+in_buf[188]*(-16)+in_buf[189]*(-6)+in_buf[190]*(-18)+in_buf[191]*(-15)+in_buf[192]*(-20)+in_buf[193]*(-31)+in_buf[194]*(-16)+in_buf[195]*(-30)+in_buf[196]*(2)+in_buf[197]*(54)+in_buf[198]*(17)+in_buf[199]*(30)+in_buf[200]*(34)+in_buf[201]*(16)+in_buf[202]*(14)+in_buf[203]*(9)+in_buf[204]*(5)+in_buf[205]*(-1)+in_buf[206]*(-14)+in_buf[207]*(0)+in_buf[208]*(0)+in_buf[209]*(10)+in_buf[210]*(7)+in_buf[211]*(9)+in_buf[212]*(-3)+in_buf[213]*(-3)+in_buf[214]*(-14)+in_buf[215]*(-17)+in_buf[216]*(-13)+in_buf[217]*(-6)+in_buf[218]*(-16)+in_buf[219]*(-22)+in_buf[220]*(-44)+in_buf[221]*(-39)+in_buf[222]*(-19)+in_buf[223]*(-40)+in_buf[224]*(5)+in_buf[225]*(34)+in_buf[226]*(36)+in_buf[227]*(38)+in_buf[228]*(27)+in_buf[229]*(8)+in_buf[230]*(0)+in_buf[231]*(3)+in_buf[232]*(3)+in_buf[233]*(-3)+in_buf[234]*(-4)+in_buf[235]*(-3)+in_buf[236]*(17)+in_buf[237]*(20)+in_buf[238]*(18)+in_buf[239]*(6)+in_buf[240]*(8)+in_buf[241]*(-12)+in_buf[242]*(-5)+in_buf[243]*(-18)+in_buf[244]*(-9)+in_buf[245]*(4)+in_buf[246]*(1)+in_buf[247]*(-60)+in_buf[248]*(-68)+in_buf[249]*(-42)+in_buf[250]*(-6)+in_buf[251]*(-9)+in_buf[252]*(7)+in_buf[253]*(37)+in_buf[254]*(45)+in_buf[255]*(16)+in_buf[256]*(11)+in_buf[257]*(9)+in_buf[258]*(3)+in_buf[259]*(6)+in_buf[260]*(-6)+in_buf[261]*(-14)+in_buf[262]*(-10)+in_buf[263]*(-6)+in_buf[264]*(10)+in_buf[265]*(13)+in_buf[266]*(15)+in_buf[267]*(-3)+in_buf[268]*(-4)+in_buf[269]*(2)+in_buf[270]*(-5)+in_buf[271]*(-1)+in_buf[272]*(20)+in_buf[273]*(11)+in_buf[274]*(2)+in_buf[275]*(-27)+in_buf[276]*(-78)+in_buf[277]*(-41)+in_buf[278]*(-30)+in_buf[279]*(-13)+in_buf[280]*(14)+in_buf[281]*(18)+in_buf[282]*(55)+in_buf[283]*(29)+in_buf[284]*(3)+in_buf[285]*(-5)+in_buf[286]*(-15)+in_buf[287]*(-11)+in_buf[288]*(-29)+in_buf[289]*(-17)+in_buf[290]*(-7)+in_buf[291]*(9)+in_buf[292]*(5)+in_buf[293]*(26)+in_buf[294]*(5)+in_buf[295]*(-23)+in_buf[296]*(-2)+in_buf[297]*(2)+in_buf[298]*(6)+in_buf[299]*(0)+in_buf[300]*(16)+in_buf[301]*(11)+in_buf[302]*(14)+in_buf[303]*(-20)+in_buf[304]*(-87)+in_buf[305]*(-47)+in_buf[306]*(-38)+in_buf[307]*(4)+in_buf[308]*(13)+in_buf[309]*(44)+in_buf[310]*(29)+in_buf[311]*(50)+in_buf[312]*(6)+in_buf[313]*(-14)+in_buf[314]*(-36)+in_buf[315]*(-34)+in_buf[316]*(-27)+in_buf[317]*(-10)+in_buf[318]*(1)+in_buf[319]*(16)+in_buf[320]*(25)+in_buf[321]*(20)+in_buf[322]*(1)+in_buf[323]*(-15)+in_buf[324]*(-11)+in_buf[325]*(6)+in_buf[326]*(6)+in_buf[327]*(2)+in_buf[328]*(6)+in_buf[329]*(4)+in_buf[330]*(-3)+in_buf[331]*(-23)+in_buf[332]*(-69)+in_buf[333]*(-74)+in_buf[334]*(-12)+in_buf[335]*(-26)+in_buf[336]*(15)+in_buf[337]*(21)+in_buf[338]*(21)+in_buf[339]*(16)+in_buf[340]*(-8)+in_buf[341]*(-10)+in_buf[342]*(-38)+in_buf[343]*(-40)+in_buf[344]*(-30)+in_buf[345]*(-9)+in_buf[346]*(7)+in_buf[347]*(22)+in_buf[348]*(25)+in_buf[349]*(15)+in_buf[350]*(7)+in_buf[351]*(15)+in_buf[352]*(9)+in_buf[353]*(19)+in_buf[354]*(13)+in_buf[355]*(-11)+in_buf[356]*(-8)+in_buf[357]*(-12)+in_buf[358]*(-4)+in_buf[359]*(-10)+in_buf[360]*(-33)+in_buf[361]*(-54)+in_buf[362]*(-25)+in_buf[363]*(-12)+in_buf[364]*(-21)+in_buf[365]*(10)+in_buf[366]*(34)+in_buf[367]*(34)+in_buf[368]*(11)+in_buf[369]*(-9)+in_buf[370]*(-23)+in_buf[371]*(-25)+in_buf[372]*(-15)+in_buf[373]*(-4)+in_buf[374]*(15)+in_buf[375]*(9)+in_buf[376]*(2)+in_buf[377]*(10)+in_buf[378]*(14)+in_buf[379]*(19)+in_buf[380]*(22)+in_buf[381]*(11)+in_buf[382]*(17)+in_buf[383]*(-1)+in_buf[384]*(-13)+in_buf[385]*(-8)+in_buf[386]*(-7)+in_buf[387]*(0)+in_buf[388]*(-23)+in_buf[389]*(-50)+in_buf[390]*(-51)+in_buf[391]*(-18)+in_buf[392]*(-10)+in_buf[393]*(11)+in_buf[394]*(6)+in_buf[395]*(21)+in_buf[396]*(9)+in_buf[397]*(2)+in_buf[398]*(-38)+in_buf[399]*(-47)+in_buf[400]*(-15)+in_buf[401]*(-2)+in_buf[402]*(8)+in_buf[403]*(13)+in_buf[404]*(9)+in_buf[405]*(12)+in_buf[406]*(10)+in_buf[407]*(25)+in_buf[408]*(2)+in_buf[409]*(3)+in_buf[410]*(15)+in_buf[411]*(11)+in_buf[412]*(0)+in_buf[413]*(0)+in_buf[414]*(-15)+in_buf[415]*(11)+in_buf[416]*(-2)+in_buf[417]*(-20)+in_buf[418]*(-41)+in_buf[419]*(-27)+in_buf[420]*(-11)+in_buf[421]*(7)+in_buf[422]*(2)+in_buf[423]*(19)+in_buf[424]*(27)+in_buf[425]*(1)+in_buf[426]*(-28)+in_buf[427]*(-34)+in_buf[428]*(-12)+in_buf[429]*(4)+in_buf[430]*(16)+in_buf[431]*(10)+in_buf[432]*(14)+in_buf[433]*(0)+in_buf[434]*(4)+in_buf[435]*(15)+in_buf[436]*(2)+in_buf[437]*(13)+in_buf[438]*(14)+in_buf[439]*(19)+in_buf[440]*(21)+in_buf[441]*(10)+in_buf[442]*(25)+in_buf[443]*(20)+in_buf[444]*(-10)+in_buf[445]*(-21)+in_buf[446]*(10)+in_buf[447]*(-33)+in_buf[448]*(8)+in_buf[449]*(23)+in_buf[450]*(20)+in_buf[451]*(24)+in_buf[452]*(30)+in_buf[453]*(-3)+in_buf[454]*(-16)+in_buf[455]*(-9)+in_buf[456]*(11)+in_buf[457]*(25)+in_buf[458]*(24)+in_buf[459]*(20)+in_buf[460]*(14)+in_buf[461]*(5)+in_buf[462]*(3)+in_buf[463]*(0)+in_buf[464]*(0)+in_buf[465]*(8)+in_buf[466]*(6)+in_buf[467]*(13)+in_buf[468]*(17)+in_buf[469]*(-9)+in_buf[470]*(-12)+in_buf[471]*(-1)+in_buf[472]*(-10)+in_buf[473]*(-50)+in_buf[474]*(-23)+in_buf[475]*(-26)+in_buf[476]*(0)+in_buf[477]*(9)+in_buf[478]*(21)+in_buf[479]*(32)+in_buf[480]*(18)+in_buf[481]*(-21)+in_buf[482]*(-31)+in_buf[483]*(-22)+in_buf[484]*(-7)+in_buf[485]*(13)+in_buf[486]*(13)+in_buf[487]*(27)+in_buf[488]*(24)+in_buf[489]*(5)+in_buf[490]*(-20)+in_buf[491]*(-7)+in_buf[492]*(6)+in_buf[493]*(13)+in_buf[494]*(-6)+in_buf[495]*(16)+in_buf[496]*(-3)+in_buf[497]*(-3)+in_buf[498]*(-5)+in_buf[499]*(0)+in_buf[500]*(-39)+in_buf[501]*(-67)+in_buf[502]*(-25)+in_buf[503]*(8)+in_buf[504]*(29)+in_buf[505]*(3)+in_buf[506]*(26)+in_buf[507]*(9)+in_buf[508]*(-11)+in_buf[509]*(-20)+in_buf[510]*(-28)+in_buf[511]*(-32)+in_buf[512]*(-14)+in_buf[513]*(-2)+in_buf[514]*(4)+in_buf[515]*(19)+in_buf[516]*(20)+in_buf[517]*(-11)+in_buf[518]*(-28)+in_buf[519]*(0)+in_buf[520]*(16)+in_buf[521]*(7)+in_buf[522]*(-4)+in_buf[523]*(5)+in_buf[524]*(-5)+in_buf[525]*(5)+in_buf[526]*(-7)+in_buf[527]*(-19)+in_buf[528]*(-63)+in_buf[529]*(-71)+in_buf[530]*(0)+in_buf[531]*(-5)+in_buf[532]*(-27)+in_buf[533]*(53)+in_buf[534]*(9)+in_buf[535]*(-1)+in_buf[536]*(0)+in_buf[537]*(-13)+in_buf[538]*(-16)+in_buf[539]*(-21)+in_buf[540]*(-11)+in_buf[541]*(0)+in_buf[542]*(5)+in_buf[543]*(0)+in_buf[544]*(1)+in_buf[545]*(-15)+in_buf[546]*(2)+in_buf[547]*(0)+in_buf[548]*(5)+in_buf[549]*(3)+in_buf[550]*(-4)+in_buf[551]*(-10)+in_buf[552]*(-1)+in_buf[553]*(7)+in_buf[554]*(-4)+in_buf[555]*(-43)+in_buf[556]*(-51)+in_buf[557]*(-50)+in_buf[558]*(-12)+in_buf[559]*(1)+in_buf[560]*(-1)+in_buf[561]*(32)+in_buf[562]*(-6)+in_buf[563]*(-6)+in_buf[564]*(-6)+in_buf[565]*(-28)+in_buf[566]*(-22)+in_buf[567]*(8)+in_buf[568]*(0)+in_buf[569]*(-2)+in_buf[570]*(-3)+in_buf[571]*(-8)+in_buf[572]*(-12)+in_buf[573]*(5)+in_buf[574]*(18)+in_buf[575]*(3)+in_buf[576]*(-7)+in_buf[577]*(-15)+in_buf[578]*(-7)+in_buf[579]*(-6)+in_buf[580]*(5)+in_buf[581]*(6)+in_buf[582]*(-8)+in_buf[583]*(-32)+in_buf[584]*(-46)+in_buf[585]*(-31)+in_buf[586]*(-10)+in_buf[587]*(-3)+in_buf[588]*(-23)+in_buf[589]*(0)+in_buf[590]*(-6)+in_buf[591]*(-6)+in_buf[592]*(-25)+in_buf[593]*(-37)+in_buf[594]*(-19)+in_buf[595]*(10)+in_buf[596]*(0)+in_buf[597]*(-26)+in_buf[598]*(-22)+in_buf[599]*(-5)+in_buf[600]*(-2)+in_buf[601]*(9)+in_buf[602]*(-4)+in_buf[603]*(-2)+in_buf[604]*(5)+in_buf[605]*(3)+in_buf[606]*(-11)+in_buf[607]*(6)+in_buf[608]*(-6)+in_buf[609]*(-10)+in_buf[610]*(-5)+in_buf[611]*(-26)+in_buf[612]*(-55)+in_buf[613]*(-37)+in_buf[614]*(16)+in_buf[615]*(5)+in_buf[616]*(-18)+in_buf[617]*(6)+in_buf[618]*(-4)+in_buf[619]*(-3)+in_buf[620]*(-3)+in_buf[621]*(-31)+in_buf[622]*(-7)+in_buf[623]*(-3)+in_buf[624]*(-11)+in_buf[625]*(-18)+in_buf[626]*(-15)+in_buf[627]*(0)+in_buf[628]*(7)+in_buf[629]*(-3)+in_buf[630]*(2)+in_buf[631]*(12)+in_buf[632]*(6)+in_buf[633]*(-3)+in_buf[634]*(-2)+in_buf[635]*(7)+in_buf[636]*(-17)+in_buf[637]*(-1)+in_buf[638]*(12)+in_buf[639]*(-8)+in_buf[640]*(-48)+in_buf[641]*(-23)+in_buf[642]*(20)+in_buf[643]*(2)+in_buf[644]*(0)+in_buf[645]*(0)+in_buf[646]*(37)+in_buf[647]*(-5)+in_buf[648]*(4)+in_buf[649]*(-3)+in_buf[650]*(-9)+in_buf[651]*(16)+in_buf[652]*(-6)+in_buf[653]*(-10)+in_buf[654]*(-1)+in_buf[655]*(0)+in_buf[656]*(-11)+in_buf[657]*(4)+in_buf[658]*(5)+in_buf[659]*(6)+in_buf[660]*(-1)+in_buf[661]*(2)+in_buf[662]*(11)+in_buf[663]*(0)+in_buf[664]*(-5)+in_buf[665]*(-17)+in_buf[666]*(-32)+in_buf[667]*(-25)+in_buf[668]*(-23)+in_buf[669]*(-9)+in_buf[670]*(-18)+in_buf[671]*(0)+in_buf[672]*(-2)+in_buf[673]*(0)+in_buf[674]*(12)+in_buf[675]*(16)+in_buf[676]*(22)+in_buf[677]*(34)+in_buf[678]*(18)+in_buf[679]*(13)+in_buf[680]*(15)+in_buf[681]*(1)+in_buf[682]*(-1)+in_buf[683]*(12)+in_buf[684]*(12)+in_buf[685]*(28)+in_buf[686]*(30)+in_buf[687]*(32)+in_buf[688]*(38)+in_buf[689]*(3)+in_buf[690]*(-19)+in_buf[691]*(-27)+in_buf[692]*(-13)+in_buf[693]*(-40)+in_buf[694]*(-41)+in_buf[695]*(-23)+in_buf[696]*(-45)+in_buf[697]*(-34)+in_buf[698]*(-28)+in_buf[699]*(-3)+in_buf[700]*(0)+in_buf[701]*(-4)+in_buf[702]*(23)+in_buf[703]*(-7)+in_buf[704]*(-4)+in_buf[705]*(18)+in_buf[706]*(7)+in_buf[707]*(12)+in_buf[708]*(13)+in_buf[709]*(9)+in_buf[710]*(37)+in_buf[711]*(29)+in_buf[712]*(0)+in_buf[713]*(3)+in_buf[714]*(-11)+in_buf[715]*(0)+in_buf[716]*(-3)+in_buf[717]*(-32)+in_buf[718]*(-7)+in_buf[719]*(11)+in_buf[720]*(-13)+in_buf[721]*(-29)+in_buf[722]*(-33)+in_buf[723]*(-10)+in_buf[724]*(-8)+in_buf[725]*(-20)+in_buf[726]*(-15)+in_buf[727]*(-3)+in_buf[728]*(0)+in_buf[729]*(0)+in_buf[730]*(2)+in_buf[731]*(3)+in_buf[732]*(-20)+in_buf[733]*(-7)+in_buf[734]*(12)+in_buf[735]*(22)+in_buf[736]*(26)+in_buf[737]*(3)+in_buf[738]*(22)+in_buf[739]*(48)+in_buf[740]*(25)+in_buf[741]*(32)+in_buf[742]*(15)+in_buf[743]*(-4)+in_buf[744]*(-1)+in_buf[745]*(-1)+in_buf[746]*(-9)+in_buf[747]*(-8)+in_buf[748]*(-1)+in_buf[749]*(-8)+in_buf[750]*(-2)+in_buf[751]*(12)+in_buf[752]*(6)+in_buf[753]*(2)+in_buf[754]*(0)+in_buf[755]*(2)+in_buf[756]*(4)+in_buf[757]*(3)+in_buf[758]*(2)+in_buf[759]*(-3)+in_buf[760]*(19)+in_buf[761]*(27)+in_buf[762]*(-9)+in_buf[763]*(-11)+in_buf[764]*(-9)+in_buf[765]*(0)+in_buf[766]*(10)+in_buf[767]*(-11)+in_buf[768]*(-8)+in_buf[769]*(14)+in_buf[770]*(-19)+in_buf[771]*(-20)+in_buf[772]*(12)+in_buf[773]*(37)+in_buf[774]*(18)+in_buf[775]*(-10)+in_buf[776]*(2)+in_buf[777]*(12)+in_buf[778]*(17)+in_buf[779]*(2)+in_buf[780]*(-3)+in_buf[781]*(-2)+in_buf[782]*(-3)+in_buf[783]*(4);
assign in_buf_weight059=in_buf[0]*(0)+in_buf[1]*(-1)+in_buf[2]*(0)+in_buf[3]*(2)+in_buf[4]*(4)+in_buf[5]*(0)+in_buf[6]*(-3)+in_buf[7]*(-2)+in_buf[8]*(-2)+in_buf[9]*(-3)+in_buf[10]*(-3)+in_buf[11]*(1)+in_buf[12]*(-11)+in_buf[13]*(-10)+in_buf[14]*(-10)+in_buf[15]*(-4)+in_buf[16]*(4)+in_buf[17]*(2)+in_buf[18]*(-3)+in_buf[19]*(-3)+in_buf[20]*(0)+in_buf[21]*(4)+in_buf[22]*(3)+in_buf[23]*(0)+in_buf[24]*(2)+in_buf[25]*(3)+in_buf[26]*(0)+in_buf[27]*(2)+in_buf[28]*(2)+in_buf[29]*(1)+in_buf[30]*(-1)+in_buf[31]*(-1)+in_buf[32]*(-8)+in_buf[33]*(0)+in_buf[34]*(-5)+in_buf[35]*(-6)+in_buf[36]*(-11)+in_buf[37]*(-13)+in_buf[38]*(-11)+in_buf[39]*(-23)+in_buf[40]*(-27)+in_buf[41]*(-3)+in_buf[42]*(17)+in_buf[43]*(-34)+in_buf[44]*(-33)+in_buf[45]*(-36)+in_buf[46]*(-16)+in_buf[47]*(-25)+in_buf[48]*(-16)+in_buf[49]*(-14)+in_buf[50]*(-10)+in_buf[51]*(-7)+in_buf[52]*(3)+in_buf[53]*(0)+in_buf[54]*(4)+in_buf[55]*(0)+in_buf[56]*(3)+in_buf[57]*(0)+in_buf[58]*(-7)+in_buf[59]*(-32)+in_buf[60]*(-32)+in_buf[61]*(-2)+in_buf[62]*(-11)+in_buf[63]*(-5)+in_buf[64]*(-9)+in_buf[65]*(-9)+in_buf[66]*(-26)+in_buf[67]*(-43)+in_buf[68]*(-20)+in_buf[69]*(-4)+in_buf[70]*(-12)+in_buf[71]*(-20)+in_buf[72]*(0)+in_buf[73]*(-5)+in_buf[74]*(-28)+in_buf[75]*(6)+in_buf[76]*(7)+in_buf[77]*(15)+in_buf[78]*(22)+in_buf[79]*(-11)+in_buf[80]*(-5)+in_buf[81]*(-3)+in_buf[82]*(-3)+in_buf[83]*(2)+in_buf[84]*(0)+in_buf[85]*(0)+in_buf[86]*(-17)+in_buf[87]*(-36)+in_buf[88]*(-25)+in_buf[89]*(-15)+in_buf[90]*(-33)+in_buf[91]*(-14)+in_buf[92]*(-45)+in_buf[93]*(-42)+in_buf[94]*(-32)+in_buf[95]*(0)+in_buf[96]*(-2)+in_buf[97]*(5)+in_buf[98]*(14)+in_buf[99]*(-21)+in_buf[100]*(-28)+in_buf[101]*(-37)+in_buf[102]*(-42)+in_buf[103]*(-30)+in_buf[104]*(-22)+in_buf[105]*(-4)+in_buf[106]*(5)+in_buf[107]*(0)+in_buf[108]*(-9)+in_buf[109]*(25)+in_buf[110]*(4)+in_buf[111]*(-1)+in_buf[112]*(-2)+in_buf[113]*(-1)+in_buf[114]*(-12)+in_buf[115]*(-2)+in_buf[116]*(-3)+in_buf[117]*(31)+in_buf[118]*(27)+in_buf[119]*(0)+in_buf[120]*(-8)+in_buf[121]*(2)+in_buf[122]*(-3)+in_buf[123]*(-14)+in_buf[124]*(10)+in_buf[125]*(20)+in_buf[126]*(1)+in_buf[127]*(-3)+in_buf[128]*(-6)+in_buf[129]*(0)+in_buf[130]*(0)+in_buf[131]*(-4)+in_buf[132]*(10)+in_buf[133]*(12)+in_buf[134]*(29)+in_buf[135]*(18)+in_buf[136]*(0)+in_buf[137]*(0)+in_buf[138]*(-23)+in_buf[139]*(-3)+in_buf[140]*(1)+in_buf[141]*(3)+in_buf[142]*(-30)+in_buf[143]*(-1)+in_buf[144]*(-18)+in_buf[145]*(21)+in_buf[146]*(25)+in_buf[147]*(-3)+in_buf[148]*(15)+in_buf[149]*(15)+in_buf[150]*(7)+in_buf[151]*(-10)+in_buf[152]*(0)+in_buf[153]*(-4)+in_buf[154]*(-5)+in_buf[155]*(2)+in_buf[156]*(-1)+in_buf[157]*(-10)+in_buf[158]*(4)+in_buf[159]*(2)+in_buf[160]*(-22)+in_buf[161]*(-13)+in_buf[162]*(-5)+in_buf[163]*(0)+in_buf[164]*(-3)+in_buf[165]*(-25)+in_buf[166]*(-23)+in_buf[167]*(-7)+in_buf[168]*(2)+in_buf[169]*(-9)+in_buf[170]*(34)+in_buf[171]*(25)+in_buf[172]*(28)+in_buf[173]*(45)+in_buf[174]*(15)+in_buf[175]*(-5)+in_buf[176]*(13)+in_buf[177]*(9)+in_buf[178]*(-7)+in_buf[179]*(-12)+in_buf[180]*(-3)+in_buf[181]*(-7)+in_buf[182]*(-23)+in_buf[183]*(-21)+in_buf[184]*(-9)+in_buf[185]*(0)+in_buf[186]*(-13)+in_buf[187]*(-13)+in_buf[188]*(-13)+in_buf[189]*(-5)+in_buf[190]*(-13)+in_buf[191]*(2)+in_buf[192]*(-13)+in_buf[193]*(-34)+in_buf[194]*(-27)+in_buf[195]*(-22)+in_buf[196]*(11)+in_buf[197]*(-26)+in_buf[198]*(28)+in_buf[199]*(38)+in_buf[200]*(18)+in_buf[201]*(28)+in_buf[202]*(16)+in_buf[203]*(5)+in_buf[204]*(3)+in_buf[205]*(9)+in_buf[206]*(0)+in_buf[207]*(0)+in_buf[208]*(-6)+in_buf[209]*(-12)+in_buf[210]*(-17)+in_buf[211]*(-12)+in_buf[212]*(-5)+in_buf[213]*(16)+in_buf[214]*(6)+in_buf[215]*(-15)+in_buf[216]*(-8)+in_buf[217]*(-2)+in_buf[218]*(4)+in_buf[219]*(3)+in_buf[220]*(-12)+in_buf[221]*(-5)+in_buf[222]*(14)+in_buf[223]*(-14)+in_buf[224]*(-4)+in_buf[225]*(19)+in_buf[226]*(17)+in_buf[227]*(4)+in_buf[228]*(9)+in_buf[229]*(25)+in_buf[230]*(12)+in_buf[231]*(-5)+in_buf[232]*(6)+in_buf[233]*(26)+in_buf[234]*(13)+in_buf[235]*(12)+in_buf[236]*(-4)+in_buf[237]*(-15)+in_buf[238]*(-19)+in_buf[239]*(0)+in_buf[240]*(2)+in_buf[241]*(3)+in_buf[242]*(-2)+in_buf[243]*(-33)+in_buf[244]*(-10)+in_buf[245]*(1)+in_buf[246]*(-16)+in_buf[247]*(0)+in_buf[248]*(7)+in_buf[249]*(4)+in_buf[250]*(3)+in_buf[251]*(-9)+in_buf[252]*(18)+in_buf[253]*(11)+in_buf[254]*(4)+in_buf[255]*(9)+in_buf[256]*(29)+in_buf[257]*(25)+in_buf[258]*(-4)+in_buf[259]*(10)+in_buf[260]*(8)+in_buf[261]*(9)+in_buf[262]*(14)+in_buf[263]*(3)+in_buf[264]*(4)+in_buf[265]*(-11)+in_buf[266]*(-21)+in_buf[267]*(4)+in_buf[268]*(5)+in_buf[269]*(20)+in_buf[270]*(0)+in_buf[271]*(-11)+in_buf[272]*(6)+in_buf[273]*(6)+in_buf[274]*(1)+in_buf[275]*(5)+in_buf[276]*(-11)+in_buf[277]*(-25)+in_buf[278]*(-3)+in_buf[279]*(-6)+in_buf[280]*(24)+in_buf[281]*(17)+in_buf[282]*(22)+in_buf[283]*(3)+in_buf[284]*(17)+in_buf[285]*(2)+in_buf[286]*(-9)+in_buf[287]*(0)+in_buf[288]*(-5)+in_buf[289]*(-2)+in_buf[290]*(-9)+in_buf[291]*(8)+in_buf[292]*(9)+in_buf[293]*(-18)+in_buf[294]*(-31)+in_buf[295]*(-6)+in_buf[296]*(8)+in_buf[297]*(23)+in_buf[298]*(2)+in_buf[299]*(2)+in_buf[300]*(8)+in_buf[301]*(18)+in_buf[302]*(9)+in_buf[303]*(-10)+in_buf[304]*(-36)+in_buf[305]*(-12)+in_buf[306]*(-30)+in_buf[307]*(-3)+in_buf[308]*(24)+in_buf[309]*(34)+in_buf[310]*(9)+in_buf[311]*(14)+in_buf[312]*(-20)+in_buf[313]*(1)+in_buf[314]*(2)+in_buf[315]*(5)+in_buf[316]*(0)+in_buf[317]*(-2)+in_buf[318]*(2)+in_buf[319]*(6)+in_buf[320]*(17)+in_buf[321]*(-21)+in_buf[322]*(-36)+in_buf[323]*(-16)+in_buf[324]*(5)+in_buf[325]*(15)+in_buf[326]*(6)+in_buf[327]*(13)+in_buf[328]*(9)+in_buf[329]*(15)+in_buf[330]*(13)+in_buf[331]*(-12)+in_buf[332]*(-60)+in_buf[333]*(-58)+in_buf[334]*(-38)+in_buf[335]*(-9)+in_buf[336]*(18)+in_buf[337]*(20)+in_buf[338]*(-2)+in_buf[339]*(7)+in_buf[340]*(-24)+in_buf[341]*(-10)+in_buf[342]*(-5)+in_buf[343]*(-5)+in_buf[344]*(1)+in_buf[345]*(-4)+in_buf[346]*(12)+in_buf[347]*(29)+in_buf[348]*(28)+in_buf[349]*(-2)+in_buf[350]*(-35)+in_buf[351]*(-21)+in_buf[352]*(4)+in_buf[353]*(11)+in_buf[354]*(10)+in_buf[355]*(8)+in_buf[356]*(15)+in_buf[357]*(19)+in_buf[358]*(24)+in_buf[359]*(-9)+in_buf[360]*(-24)+in_buf[361]*(-23)+in_buf[362]*(-17)+in_buf[363]*(-7)+in_buf[364]*(3)+in_buf[365]*(13)+in_buf[366]*(24)+in_buf[367]*(-4)+in_buf[368]*(-1)+in_buf[369]*(-1)+in_buf[370]*(-2)+in_buf[371]*(-2)+in_buf[372]*(3)+in_buf[373]*(11)+in_buf[374]*(21)+in_buf[375]*(21)+in_buf[376]*(6)+in_buf[377]*(-30)+in_buf[378]*(-49)+in_buf[379]*(-38)+in_buf[380]*(1)+in_buf[381]*(25)+in_buf[382]*(19)+in_buf[383]*(9)+in_buf[384]*(21)+in_buf[385]*(25)+in_buf[386]*(2)+in_buf[387]*(-28)+in_buf[388]*(-16)+in_buf[389]*(-20)+in_buf[390]*(-18)+in_buf[391]*(-9)+in_buf[392]*(-9)+in_buf[393]*(16)+in_buf[394]*(26)+in_buf[395]*(-8)+in_buf[396]*(8)+in_buf[397]*(3)+in_buf[398]*(-13)+in_buf[399]*(17)+in_buf[400]*(24)+in_buf[401]*(22)+in_buf[402]*(21)+in_buf[403]*(10)+in_buf[404]*(1)+in_buf[405]*(-21)+in_buf[406]*(-37)+in_buf[407]*(-29)+in_buf[408]*(3)+in_buf[409]*(25)+in_buf[410]*(21)+in_buf[411]*(34)+in_buf[412]*(27)+in_buf[413]*(9)+in_buf[414]*(-20)+in_buf[415]*(-36)+in_buf[416]*(-28)+in_buf[417]*(-30)+in_buf[418]*(-27)+in_buf[419]*(-10)+in_buf[420]*(-10)+in_buf[421]*(-7)+in_buf[422]*(21)+in_buf[423]*(7)+in_buf[424]*(-16)+in_buf[425]*(-12)+in_buf[426]*(-9)+in_buf[427]*(19)+in_buf[428]*(11)+in_buf[429]*(22)+in_buf[430]*(23)+in_buf[431]*(7)+in_buf[432]*(-6)+in_buf[433]*(-10)+in_buf[434]*(-36)+in_buf[435]*(-12)+in_buf[436]*(16)+in_buf[437]*(30)+in_buf[438]*(26)+in_buf[439]*(34)+in_buf[440]*(20)+in_buf[441]*(4)+in_buf[442]*(-3)+in_buf[443]*(-39)+in_buf[444]*(-43)+in_buf[445]*(-30)+in_buf[446]*(11)+in_buf[447]*(-29)+in_buf[448]*(19)+in_buf[449]*(-8)+in_buf[450]*(12)+in_buf[451]*(-7)+in_buf[452]*(-8)+in_buf[453]*(-5)+in_buf[454]*(7)+in_buf[455]*(29)+in_buf[456]*(22)+in_buf[457]*(21)+in_buf[458]*(9)+in_buf[459]*(0)+in_buf[460]*(-11)+in_buf[461]*(-40)+in_buf[462]*(-25)+in_buf[463]*(15)+in_buf[464]*(21)+in_buf[465]*(31)+in_buf[466]*(29)+in_buf[467]*(33)+in_buf[468]*(28)+in_buf[469]*(14)+in_buf[470]*(2)+in_buf[471]*(-12)+in_buf[472]*(-15)+in_buf[473]*(-19)+in_buf[474]*(-17)+in_buf[475]*(-28)+in_buf[476]*(3)+in_buf[477]*(-11)+in_buf[478]*(34)+in_buf[479]*(-27)+in_buf[480]*(4)+in_buf[481]*(-12)+in_buf[482]*(-11)+in_buf[483]*(4)+in_buf[484]*(21)+in_buf[485]*(26)+in_buf[486]*(18)+in_buf[487]*(-15)+in_buf[488]*(-47)+in_buf[489]*(-51)+in_buf[490]*(-12)+in_buf[491]*(21)+in_buf[492]*(25)+in_buf[493]*(27)+in_buf[494]*(39)+in_buf[495]*(15)+in_buf[496]*(7)+in_buf[497]*(6)+in_buf[498]*(6)+in_buf[499]*(-8)+in_buf[500]*(1)+in_buf[501]*(-6)+in_buf[502]*(-7)+in_buf[503]*(-26)+in_buf[504]*(0)+in_buf[505]*(-5)+in_buf[506]*(22)+in_buf[507]*(-15)+in_buf[508]*(-5)+in_buf[509]*(-19)+in_buf[510]*(-24)+in_buf[511]*(-3)+in_buf[512]*(1)+in_buf[513]*(5)+in_buf[514]*(-17)+in_buf[515]*(-44)+in_buf[516]*(-64)+in_buf[517]*(-39)+in_buf[518]*(4)+in_buf[519]*(21)+in_buf[520]*(33)+in_buf[521]*(27)+in_buf[522]*(26)+in_buf[523]*(9)+in_buf[524]*(-8)+in_buf[525]*(8)+in_buf[526]*(-3)+in_buf[527]*(-19)+in_buf[528]*(-10)+in_buf[529]*(-48)+in_buf[530]*(-14)+in_buf[531]*(3)+in_buf[532]*(0)+in_buf[533]*(30)+in_buf[534]*(13)+in_buf[535]*(22)+in_buf[536]*(-3)+in_buf[537]*(-11)+in_buf[538]*(-5)+in_buf[539]*(5)+in_buf[540]*(6)+in_buf[541]*(-7)+in_buf[542]*(-29)+in_buf[543]*(-44)+in_buf[544]*(-73)+in_buf[545]*(-38)+in_buf[546]*(7)+in_buf[547]*(23)+in_buf[548]*(20)+in_buf[549]*(16)+in_buf[550]*(1)+in_buf[551]*(-2)+in_buf[552]*(-20)+in_buf[553]*(-5)+in_buf[554]*(-32)+in_buf[555]*(-50)+in_buf[556]*(-18)+in_buf[557]*(-43)+in_buf[558]*(-7)+in_buf[559]*(-5)+in_buf[560]*(-1)+in_buf[561]*(1)+in_buf[562]*(31)+in_buf[563]*(6)+in_buf[564]*(-14)+in_buf[565]*(-5)+in_buf[566]*(-9)+in_buf[567]*(-2)+in_buf[568]*(-14)+in_buf[569]*(-18)+in_buf[570]*(-19)+in_buf[571]*(-25)+in_buf[572]*(-16)+in_buf[573]*(-7)+in_buf[574]*(11)+in_buf[575]*(10)+in_buf[576]*(21)+in_buf[577]*(15)+in_buf[578]*(9)+in_buf[579]*(-5)+in_buf[580]*(-24)+in_buf[581]*(-26)+in_buf[582]*(-31)+in_buf[583]*(-35)+in_buf[584]*(0)+in_buf[585]*(-31)+in_buf[586]*(12)+in_buf[587]*(-3)+in_buf[588]*(-5)+in_buf[589]*(9)+in_buf[590]*(3)+in_buf[591]*(-1)+in_buf[592]*(-1)+in_buf[593]*(7)+in_buf[594]*(-18)+in_buf[595]*(-29)+in_buf[596]*(-13)+in_buf[597]*(-24)+in_buf[598]*(-3)+in_buf[599]*(3)+in_buf[600]*(0)+in_buf[601]*(14)+in_buf[602]*(10)+in_buf[603]*(0)+in_buf[604]*(16)+in_buf[605]*(3)+in_buf[606]*(-6)+in_buf[607]*(-1)+in_buf[608]*(-18)+in_buf[609]*(-7)+in_buf[610]*(2)+in_buf[611]*(-7)+in_buf[612]*(3)+in_buf[613]*(-7)+in_buf[614]*(-28)+in_buf[615]*(0)+in_buf[616]*(-3)+in_buf[617]*(-19)+in_buf[618]*(5)+in_buf[619]*(-2)+in_buf[620]*(-9)+in_buf[621]*(-8)+in_buf[622]*(-4)+in_buf[623]*(-12)+in_buf[624]*(-16)+in_buf[625]*(-19)+in_buf[626]*(-8)+in_buf[627]*(5)+in_buf[628]*(13)+in_buf[629]*(23)+in_buf[630]*(12)+in_buf[631]*(9)+in_buf[632]*(7)+in_buf[633]*(-4)+in_buf[634]*(-9)+in_buf[635]*(0)+in_buf[636]*(-6)+in_buf[637]*(-2)+in_buf[638]*(6)+in_buf[639]*(-23)+in_buf[640]*(6)+in_buf[641]*(-4)+in_buf[642]*(0)+in_buf[643]*(4)+in_buf[644]*(1)+in_buf[645]*(-1)+in_buf[646]*(-29)+in_buf[647]*(-3)+in_buf[648]*(-26)+in_buf[649]*(2)+in_buf[650]*(11)+in_buf[651]*(5)+in_buf[652]*(-2)+in_buf[653]*(-8)+in_buf[654]*(-6)+in_buf[655]*(5)+in_buf[656]*(24)+in_buf[657]*(17)+in_buf[658]*(18)+in_buf[659]*(7)+in_buf[660]*(7)+in_buf[661]*(0)+in_buf[662]*(-4)+in_buf[663]*(11)+in_buf[664]*(0)+in_buf[665]*(10)+in_buf[666]*(-22)+in_buf[667]*(-20)+in_buf[668]*(-3)+in_buf[669]*(-3)+in_buf[670]*(-9)+in_buf[671]*(-2)+in_buf[672]*(-1)+in_buf[673]*(-3)+in_buf[674]*(11)+in_buf[675]*(-3)+in_buf[676]*(3)+in_buf[677]*(1)+in_buf[678]*(-13)+in_buf[679]*(-23)+in_buf[680]*(-16)+in_buf[681]*(12)+in_buf[682]*(5)+in_buf[683]*(1)+in_buf[684]*(9)+in_buf[685]*(6)+in_buf[686]*(-11)+in_buf[687]*(-13)+in_buf[688]*(15)+in_buf[689]*(11)+in_buf[690]*(0)+in_buf[691]*(12)+in_buf[692]*(19)+in_buf[693]*(31)+in_buf[694]*(-7)+in_buf[695]*(-27)+in_buf[696]*(0)+in_buf[697]*(18)+in_buf[698]*(9)+in_buf[699]*(4)+in_buf[700]*(0)+in_buf[701]*(-2)+in_buf[702]*(-8)+in_buf[703]*(-13)+in_buf[704]*(-1)+in_buf[705]*(-13)+in_buf[706]*(-24)+in_buf[707]*(-54)+in_buf[708]*(-12)+in_buf[709]*(-7)+in_buf[710]*(-14)+in_buf[711]*(0)+in_buf[712]*(-8)+in_buf[713]*(-4)+in_buf[714]*(19)+in_buf[715]*(10)+in_buf[716]*(6)+in_buf[717]*(12)+in_buf[718]*(9)+in_buf[719]*(-30)+in_buf[720]*(-24)+in_buf[721]*(-23)+in_buf[722]*(-22)+in_buf[723]*(-30)+in_buf[724]*(-45)+in_buf[725]*(5)+in_buf[726]*(16)+in_buf[727]*(-2)+in_buf[728]*(2)+in_buf[729]*(0)+in_buf[730]*(1)+in_buf[731]*(2)+in_buf[732]*(-2)+in_buf[733]*(-25)+in_buf[734]*(-11)+in_buf[735]*(3)+in_buf[736]*(-11)+in_buf[737]*(-12)+in_buf[738]*(-17)+in_buf[739]*(-27)+in_buf[740]*(-33)+in_buf[741]*(-35)+in_buf[742]*(-35)+in_buf[743]*(-19)+in_buf[744]*(-16)+in_buf[745]*(-30)+in_buf[746]*(-20)+in_buf[747]*(-16)+in_buf[748]*(-16)+in_buf[749]*(-23)+in_buf[750]*(-39)+in_buf[751]*(-40)+in_buf[752]*(-10)+in_buf[753]*(4)+in_buf[754]*(3)+in_buf[755]*(1)+in_buf[756]*(0)+in_buf[757]*(-1)+in_buf[758]*(0)+in_buf[759]*(-2)+in_buf[760]*(8)+in_buf[761]*(29)+in_buf[762]*(-3)+in_buf[763]*(-16)+in_buf[764]*(-18)+in_buf[765]*(6)+in_buf[766]*(-10)+in_buf[767]*(-16)+in_buf[768]*(-19)+in_buf[769]*(-1)+in_buf[770]*(-35)+in_buf[771]*(-35)+in_buf[772]*(-17)+in_buf[773]*(23)+in_buf[774]*(28)+in_buf[775]*(3)+in_buf[776]*(19)+in_buf[777]*(27)+in_buf[778]*(10)+in_buf[779]*(32)+in_buf[780]*(4)+in_buf[781]*(0)+in_buf[782]*(2)+in_buf[783]*(4);
assign in_buf_weight060=in_buf[0]*(2)+in_buf[1]*(1)+in_buf[2]*(3)+in_buf[3]*(-1)+in_buf[4]*(1)+in_buf[5]*(-1)+in_buf[6]*(0)+in_buf[7]*(3)+in_buf[8]*(4)+in_buf[9]*(-1)+in_buf[10]*(1)+in_buf[11]*(-1)+in_buf[12]*(-9)+in_buf[13]*(-6)+in_buf[14]*(12)+in_buf[15]*(3)+in_buf[16]*(2)+in_buf[17]*(-3)+in_buf[18]*(0)+in_buf[19]*(4)+in_buf[20]*(1)+in_buf[21]*(0)+in_buf[22]*(1)+in_buf[23]*(3)+in_buf[24]*(-2)+in_buf[25]*(5)+in_buf[26]*(-1)+in_buf[27]*(2)+in_buf[28]*(0)+in_buf[29]*(4)+in_buf[30]*(1)+in_buf[31]*(4)+in_buf[32]*(6)+in_buf[33]*(-7)+in_buf[34]*(-9)+in_buf[35]*(-8)+in_buf[36]*(-8)+in_buf[37]*(0)+in_buf[38]*(16)+in_buf[39]*(4)+in_buf[40]*(5)+in_buf[41]*(13)+in_buf[42]*(10)+in_buf[43]*(-13)+in_buf[44]*(-15)+in_buf[45]*(-11)+in_buf[46]*(-6)+in_buf[47]*(-13)+in_buf[48]*(-16)+in_buf[49]*(-19)+in_buf[50]*(-11)+in_buf[51]*(-15)+in_buf[52]*(2)+in_buf[53]*(-3)+in_buf[54]*(-2)+in_buf[55]*(3)+in_buf[56]*(-2)+in_buf[57]*(2)+in_buf[58]*(0)+in_buf[59]*(-14)+in_buf[60]*(-10)+in_buf[61]*(-4)+in_buf[62]*(-9)+in_buf[63]*(-9)+in_buf[64]*(8)+in_buf[65]*(21)+in_buf[66]*(-10)+in_buf[67]*(-15)+in_buf[68]*(-16)+in_buf[69]*(-4)+in_buf[70]*(18)+in_buf[71]*(0)+in_buf[72]*(3)+in_buf[73]*(18)+in_buf[74]*(9)+in_buf[75]*(10)+in_buf[76]*(8)+in_buf[77]*(0)+in_buf[78]*(-23)+in_buf[79]*(-40)+in_buf[80]*(-3)+in_buf[81]*(-3)+in_buf[82]*(-1)+in_buf[83]*(-1)+in_buf[84]*(-3)+in_buf[85]*(0)+in_buf[86]*(-22)+in_buf[87]*(-17)+in_buf[88]*(17)+in_buf[89]*(5)+in_buf[90]*(-17)+in_buf[91]*(6)+in_buf[92]*(-7)+in_buf[93]*(15)+in_buf[94]*(5)+in_buf[95]*(11)+in_buf[96]*(-1)+in_buf[97]*(12)+in_buf[98]*(12)+in_buf[99]*(10)+in_buf[100]*(19)+in_buf[101]*(4)+in_buf[102]*(-9)+in_buf[103]*(-7)+in_buf[104]*(16)+in_buf[105]*(25)+in_buf[106]*(2)+in_buf[107]*(-23)+in_buf[108]*(29)+in_buf[109]*(27)+in_buf[110]*(30)+in_buf[111]*(-1)+in_buf[112]*(-3)+in_buf[113]*(-3)+in_buf[114]*(-28)+in_buf[115]*(-25)+in_buf[116]*(-20)+in_buf[117]*(-20)+in_buf[118]*(0)+in_buf[119]*(9)+in_buf[120]*(0)+in_buf[121]*(20)+in_buf[122]*(8)+in_buf[123]*(16)+in_buf[124]*(22)+in_buf[125]*(12)+in_buf[126]*(-1)+in_buf[127]*(15)+in_buf[128]*(14)+in_buf[129]*(6)+in_buf[130]*(-22)+in_buf[131]*(-25)+in_buf[132]*(-12)+in_buf[133]*(3)+in_buf[134]*(-11)+in_buf[135]*(23)+in_buf[136]*(37)+in_buf[137]*(28)+in_buf[138]*(-14)+in_buf[139]*(15)+in_buf[140]*(3)+in_buf[141]*(4)+in_buf[142]*(-29)+in_buf[143]*(20)+in_buf[144]*(10)+in_buf[145]*(-5)+in_buf[146]*(9)+in_buf[147]*(8)+in_buf[148]*(14)+in_buf[149]*(14)+in_buf[150]*(19)+in_buf[151]*(8)+in_buf[152]*(-14)+in_buf[153]*(-47)+in_buf[154]*(-35)+in_buf[155]*(1)+in_buf[156]*(21)+in_buf[157]*(13)+in_buf[158]*(-1)+in_buf[159]*(-7)+in_buf[160]*(-1)+in_buf[161]*(9)+in_buf[162]*(5)+in_buf[163]*(29)+in_buf[164]*(28)+in_buf[165]*(32)+in_buf[166]*(17)+in_buf[167]*(21)+in_buf[168]*(0)+in_buf[169]*(4)+in_buf[170]*(19)+in_buf[171]*(15)+in_buf[172]*(44)+in_buf[173]*(48)+in_buf[174]*(19)+in_buf[175]*(13)+in_buf[176]*(12)+in_buf[177]*(6)+in_buf[178]*(-22)+in_buf[179]*(-27)+in_buf[180]*(-44)+in_buf[181]*(-68)+in_buf[182]*(-61)+in_buf[183]*(-21)+in_buf[184]*(9)+in_buf[185]*(-5)+in_buf[186]*(-6)+in_buf[187]*(-4)+in_buf[188]*(1)+in_buf[189]*(4)+in_buf[190]*(21)+in_buf[191]*(24)+in_buf[192]*(26)+in_buf[193]*(31)+in_buf[194]*(9)+in_buf[195]*(19)+in_buf[196]*(2)+in_buf[197]*(3)+in_buf[198]*(-1)+in_buf[199]*(5)+in_buf[200]*(20)+in_buf[201]*(28)+in_buf[202]*(4)+in_buf[203]*(3)+in_buf[204]*(25)+in_buf[205]*(17)+in_buf[206]*(6)+in_buf[207]*(-23)+in_buf[208]*(-37)+in_buf[209]*(-53)+in_buf[210]*(-42)+in_buf[211]*(-23)+in_buf[212]*(0)+in_buf[213]*(9)+in_buf[214]*(-1)+in_buf[215]*(-14)+in_buf[216]*(-5)+in_buf[217]*(7)+in_buf[218]*(24)+in_buf[219]*(-1)+in_buf[220]*(15)+in_buf[221]*(39)+in_buf[222]*(26)+in_buf[223]*(22)+in_buf[224]*(36)+in_buf[225]*(-18)+in_buf[226]*(-12)+in_buf[227]*(0)+in_buf[228]*(0)+in_buf[229]*(4)+in_buf[230]*(0)+in_buf[231]*(-3)+in_buf[232]*(14)+in_buf[233]*(39)+in_buf[234]*(18)+in_buf[235]*(-1)+in_buf[236]*(-24)+in_buf[237]*(-34)+in_buf[238]*(-27)+in_buf[239]*(-16)+in_buf[240]*(0)+in_buf[241]*(7)+in_buf[242]*(-11)+in_buf[243]*(-13)+in_buf[244]*(14)+in_buf[245]*(11)+in_buf[246]*(8)+in_buf[247]*(19)+in_buf[248]*(15)+in_buf[249]*(38)+in_buf[250]*(18)+in_buf[251]*(-7)+in_buf[252]*(-5)+in_buf[253]*(0)+in_buf[254]*(-20)+in_buf[255]*(3)+in_buf[256]*(-12)+in_buf[257]*(3)+in_buf[258]*(-14)+in_buf[259]*(4)+in_buf[260]*(14)+in_buf[261]*(24)+in_buf[262]*(18)+in_buf[263]*(2)+in_buf[264]*(-27)+in_buf[265]*(-24)+in_buf[266]*(-8)+in_buf[267]*(-5)+in_buf[268]*(18)+in_buf[269]*(12)+in_buf[270]*(1)+in_buf[271]*(4)+in_buf[272]*(22)+in_buf[273]*(16)+in_buf[274]*(-4)+in_buf[275]*(5)+in_buf[276]*(29)+in_buf[277]*(31)+in_buf[278]*(22)+in_buf[279]*(-14)+in_buf[280]*(-4)+in_buf[281]*(-7)+in_buf[282]*(-24)+in_buf[283]*(17)+in_buf[284]*(9)+in_buf[285]*(7)+in_buf[286]*(-4)+in_buf[287]*(12)+in_buf[288]*(31)+in_buf[289]*(28)+in_buf[290]*(16)+in_buf[291]*(-1)+in_buf[292]*(-30)+in_buf[293]*(-29)+in_buf[294]*(-11)+in_buf[295]*(14)+in_buf[296]*(22)+in_buf[297]*(16)+in_buf[298]*(1)+in_buf[299]*(3)+in_buf[300]*(9)+in_buf[301]*(10)+in_buf[302]*(-2)+in_buf[303]*(-28)+in_buf[304]*(16)+in_buf[305]*(38)+in_buf[306]*(50)+in_buf[307]*(-21)+in_buf[308]*(-5)+in_buf[309]*(27)+in_buf[310]*(-36)+in_buf[311]*(0)+in_buf[312]*(-11)+in_buf[313]*(-2)+in_buf[314]*(-14)+in_buf[315]*(-9)+in_buf[316]*(14)+in_buf[317]*(15)+in_buf[318]*(22)+in_buf[319]*(-5)+in_buf[320]*(-32)+in_buf[321]*(-39)+in_buf[322]*(-32)+in_buf[323]*(-2)+in_buf[324]*(13)+in_buf[325]*(-7)+in_buf[326]*(-20)+in_buf[327]*(-4)+in_buf[328]*(-21)+in_buf[329]*(-24)+in_buf[330]*(-37)+in_buf[331]*(-48)+in_buf[332]*(-36)+in_buf[333]*(22)+in_buf[334]*(52)+in_buf[335]*(-19)+in_buf[336]*(-3)+in_buf[337]*(4)+in_buf[338]*(-17)+in_buf[339]*(-7)+in_buf[340]*(-26)+in_buf[341]*(-17)+in_buf[342]*(-19)+in_buf[343]*(8)+in_buf[344]*(12)+in_buf[345]*(10)+in_buf[346]*(29)+in_buf[347]*(3)+in_buf[348]*(-4)+in_buf[349]*(-9)+in_buf[350]*(-28)+in_buf[351]*(-10)+in_buf[352]*(-5)+in_buf[353]*(-16)+in_buf[354]*(-22)+in_buf[355]*(-14)+in_buf[356]*(-26)+in_buf[357]*(-29)+in_buf[358]*(-28)+in_buf[359]*(-47)+in_buf[360]*(-33)+in_buf[361]*(6)+in_buf[362]*(7)+in_buf[363]*(-20)+in_buf[364]*(4)+in_buf[365]*(4)+in_buf[366]*(-2)+in_buf[367]*(0)+in_buf[368]*(-38)+in_buf[369]*(-2)+in_buf[370]*(11)+in_buf[371]*(14)+in_buf[372]*(15)+in_buf[373]*(7)+in_buf[374]*(16)+in_buf[375]*(11)+in_buf[376]*(28)+in_buf[377]*(-5)+in_buf[378]*(-24)+in_buf[379]*(-11)+in_buf[380]*(-8)+in_buf[381]*(-2)+in_buf[382]*(9)+in_buf[383]*(-13)+in_buf[384]*(-7)+in_buf[385]*(-19)+in_buf[386]*(-5)+in_buf[387]*(6)+in_buf[388]*(15)+in_buf[389]*(-5)+in_buf[390]*(6)+in_buf[391]*(16)+in_buf[392]*(1)+in_buf[393]*(3)+in_buf[394]*(1)+in_buf[395]*(19)+in_buf[396]*(-10)+in_buf[397]*(25)+in_buf[398]*(15)+in_buf[399]*(24)+in_buf[400]*(9)+in_buf[401]*(15)+in_buf[402]*(4)+in_buf[403]*(14)+in_buf[404]*(23)+in_buf[405]*(7)+in_buf[406]*(-10)+in_buf[407]*(3)+in_buf[408]*(1)+in_buf[409]*(8)+in_buf[410]*(0)+in_buf[411]*(-3)+in_buf[412]*(-3)+in_buf[413]*(-4)+in_buf[414]*(16)+in_buf[415]*(15)+in_buf[416]*(55)+in_buf[417]*(30)+in_buf[418]*(26)+in_buf[419]*(7)+in_buf[420]*(0)+in_buf[421]*(6)+in_buf[422]*(24)+in_buf[423]*(46)+in_buf[424]*(23)+in_buf[425]*(10)+in_buf[426]*(2)+in_buf[427]*(12)+in_buf[428]*(8)+in_buf[429]*(9)+in_buf[430]*(8)+in_buf[431]*(24)+in_buf[432]*(32)+in_buf[433]*(22)+in_buf[434]*(0)+in_buf[435]*(-2)+in_buf[436]*(11)+in_buf[437]*(24)+in_buf[438]*(4)+in_buf[439]*(2)+in_buf[440]*(2)+in_buf[441]*(11)+in_buf[442]*(26)+in_buf[443]*(43)+in_buf[444]*(48)+in_buf[445]*(42)+in_buf[446]*(26)+in_buf[447]*(24)+in_buf[448]*(-9)+in_buf[449]*(3)+in_buf[450]*(-5)+in_buf[451]*(37)+in_buf[452]*(9)+in_buf[453]*(0)+in_buf[454]*(-6)+in_buf[455]*(-2)+in_buf[456]*(8)+in_buf[457]*(9)+in_buf[458]*(7)+in_buf[459]*(19)+in_buf[460]*(16)+in_buf[461]*(11)+in_buf[462]*(7)+in_buf[463]*(19)+in_buf[464]*(17)+in_buf[465]*(16)+in_buf[466]*(8)+in_buf[467]*(12)+in_buf[468]*(25)+in_buf[469]*(48)+in_buf[470]*(36)+in_buf[471]*(43)+in_buf[472]*(16)+in_buf[473]*(29)+in_buf[474]*(48)+in_buf[475]*(26)+in_buf[476]*(-3)+in_buf[477]*(-3)+in_buf[478]*(25)+in_buf[479]*(9)+in_buf[480]*(16)+in_buf[481]*(5)+in_buf[482]*(7)+in_buf[483]*(7)+in_buf[484]*(3)+in_buf[485]*(10)+in_buf[486]*(2)+in_buf[487]*(-1)+in_buf[488]*(2)+in_buf[489]*(-5)+in_buf[490]*(-4)+in_buf[491]*(7)+in_buf[492]*(17)+in_buf[493]*(-3)+in_buf[494]*(14)+in_buf[495]*(-5)+in_buf[496]*(7)+in_buf[497]*(29)+in_buf[498]*(24)+in_buf[499]*(15)+in_buf[500]*(-8)+in_buf[501]*(-2)+in_buf[502]*(11)+in_buf[503]*(21)+in_buf[504]*(-31)+in_buf[505]*(-11)+in_buf[506]*(21)+in_buf[507]*(2)+in_buf[508]*(-1)+in_buf[509]*(21)+in_buf[510]*(19)+in_buf[511]*(4)+in_buf[512]*(2)+in_buf[513]*(4)+in_buf[514]*(1)+in_buf[515]*(5)+in_buf[516]*(22)+in_buf[517]*(14)+in_buf[518]*(11)+in_buf[519]*(4)+in_buf[520]*(9)+in_buf[521]*(-18)+in_buf[522]*(-5)+in_buf[523]*(-13)+in_buf[524]*(-10)+in_buf[525]*(2)+in_buf[526]*(-12)+in_buf[527]*(9)+in_buf[528]*(9)+in_buf[529]*(-6)+in_buf[530]*(-22)+in_buf[531]*(8)+in_buf[532]*(-12)+in_buf[533]*(-11)+in_buf[534]*(-22)+in_buf[535]*(23)+in_buf[536]*(5)+in_buf[537]*(11)+in_buf[538]*(4)+in_buf[539]*(-2)+in_buf[540]*(-9)+in_buf[541]*(0)+in_buf[542]*(10)+in_buf[543]*(20)+in_buf[544]*(3)+in_buf[545]*(1)+in_buf[546]*(18)+in_buf[547]*(7)+in_buf[548]*(0)+in_buf[549]*(-8)+in_buf[550]*(4)+in_buf[551]*(-20)+in_buf[552]*(-2)+in_buf[553]*(3)+in_buf[554]*(-5)+in_buf[555]*(9)+in_buf[556]*(-1)+in_buf[557]*(-1)+in_buf[558]*(31)+in_buf[559]*(2)+in_buf[560]*(4)+in_buf[561]*(20)+in_buf[562]*(3)+in_buf[563]*(26)+in_buf[564]*(-14)+in_buf[565]*(-18)+in_buf[566]*(-25)+in_buf[567]*(-12)+in_buf[568]*(-7)+in_buf[569]*(8)+in_buf[570]*(12)+in_buf[571]*(19)+in_buf[572]*(14)+in_buf[573]*(5)+in_buf[574]*(1)+in_buf[575]*(8)+in_buf[576]*(-8)+in_buf[577]*(-3)+in_buf[578]*(4)+in_buf[579]*(-16)+in_buf[580]*(0)+in_buf[581]*(7)+in_buf[582]*(0)+in_buf[583]*(0)+in_buf[584]*(-22)+in_buf[585]*(-8)+in_buf[586]*(28)+in_buf[587]*(3)+in_buf[588]*(-15)+in_buf[589]*(-8)+in_buf[590]*(1)+in_buf[591]*(23)+in_buf[592]*(6)+in_buf[593]*(-17)+in_buf[594]*(-22)+in_buf[595]*(-19)+in_buf[596]*(-26)+in_buf[597]*(0)+in_buf[598]*(4)+in_buf[599]*(17)+in_buf[600]*(18)+in_buf[601]*(10)+in_buf[602]*(0)+in_buf[603]*(-4)+in_buf[604]*(0)+in_buf[605]*(5)+in_buf[606]*(-4)+in_buf[607]*(-2)+in_buf[608]*(1)+in_buf[609]*(20)+in_buf[610]*(20)+in_buf[611]*(8)+in_buf[612]*(-13)+in_buf[613]*(11)+in_buf[614]*(32)+in_buf[615]*(3)+in_buf[616]*(-18)+in_buf[617]*(-15)+in_buf[618]*(10)+in_buf[619]*(19)+in_buf[620]*(-10)+in_buf[621]*(-38)+in_buf[622]*(-29)+in_buf[623]*(-21)+in_buf[624]*(-32)+in_buf[625]*(-22)+in_buf[626]*(-1)+in_buf[627]*(1)+in_buf[628]*(0)+in_buf[629]*(3)+in_buf[630]*(-3)+in_buf[631]*(4)+in_buf[632]*(8)+in_buf[633]*(-3)+in_buf[634]*(-16)+in_buf[635]*(-1)+in_buf[636]*(-3)+in_buf[637]*(11)+in_buf[638]*(17)+in_buf[639]*(5)+in_buf[640]*(-15)+in_buf[641]*(-3)+in_buf[642]*(34)+in_buf[643]*(0)+in_buf[644]*(-1)+in_buf[645]*(-2)+in_buf[646]*(2)+in_buf[647]*(11)+in_buf[648]*(9)+in_buf[649]*(-33)+in_buf[650]*(-22)+in_buf[651]*(-36)+in_buf[652]*(-37)+in_buf[653]*(-26)+in_buf[654]*(-12)+in_buf[655]*(-30)+in_buf[656]*(-16)+in_buf[657]*(-1)+in_buf[658]*(14)+in_buf[659]*(-7)+in_buf[660]*(-4)+in_buf[661]*(-15)+in_buf[662]*(-12)+in_buf[663]*(-16)+in_buf[664]*(-26)+in_buf[665]*(2)+in_buf[666]*(3)+in_buf[667]*(-13)+in_buf[668]*(-19)+in_buf[669]*(14)+in_buf[670]*(17)+in_buf[671]*(-1)+in_buf[672]*(-2)+in_buf[673]*(-2)+in_buf[674]*(8)+in_buf[675]*(7)+in_buf[676]*(0)+in_buf[677]*(-11)+in_buf[678]*(-33)+in_buf[679]*(-41)+in_buf[680]*(-47)+in_buf[681]*(-33)+in_buf[682]*(-48)+in_buf[683]*(-21)+in_buf[684]*(-20)+in_buf[685]*(-11)+in_buf[686]*(12)+in_buf[687]*(1)+in_buf[688]*(-2)+in_buf[689]*(0)+in_buf[690]*(0)+in_buf[691]*(-18)+in_buf[692]*(-16)+in_buf[693]*(-6)+in_buf[694]*(0)+in_buf[695]*(-21)+in_buf[696]*(12)+in_buf[697]*(10)+in_buf[698]*(15)+in_buf[699]*(-2)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(0)+in_buf[703]*(6)+in_buf[704]*(-7)+in_buf[705]*(-27)+in_buf[706]*(-37)+in_buf[707]*(-42)+in_buf[708]*(-31)+in_buf[709]*(-34)+in_buf[710]*(-56)+in_buf[711]*(-20)+in_buf[712]*(-51)+in_buf[713]*(-31)+in_buf[714]*(-5)+in_buf[715]*(8)+in_buf[716]*(-5)+in_buf[717]*(1)+in_buf[718]*(-10)+in_buf[719]*(-39)+in_buf[720]*(-33)+in_buf[721]*(-20)+in_buf[722]*(-1)+in_buf[723]*(14)+in_buf[724]*(12)+in_buf[725]*(-3)+in_buf[726]*(17)+in_buf[727]*(4)+in_buf[728]*(-3)+in_buf[729]*(-1)+in_buf[730]*(-2)+in_buf[731]*(1)+in_buf[732]*(-10)+in_buf[733]*(-26)+in_buf[734]*(-38)+in_buf[735]*(-49)+in_buf[736]*(-61)+in_buf[737]*(-63)+in_buf[738]*(-61)+in_buf[739]*(-41)+in_buf[740]*(-36)+in_buf[741]*(-54)+in_buf[742]*(-79)+in_buf[743]*(-54)+in_buf[744]*(-26)+in_buf[745]*(-18)+in_buf[746]*(-42)+in_buf[747]*(-56)+in_buf[748]*(-49)+in_buf[749]*(-38)+in_buf[750]*(-36)+in_buf[751]*(-2)+in_buf[752]*(-20)+in_buf[753]*(0)+in_buf[754]*(4)+in_buf[755]*(0)+in_buf[756]*(4)+in_buf[757]*(3)+in_buf[758]*(0)+in_buf[759]*(4)+in_buf[760]*(-3)+in_buf[761]*(2)+in_buf[762]*(-13)+in_buf[763]*(-12)+in_buf[764]*(-14)+in_buf[765]*(-14)+in_buf[766]*(-33)+in_buf[767]*(-29)+in_buf[768]*(-16)+in_buf[769]*(-25)+in_buf[770]*(-58)+in_buf[771]*(-43)+in_buf[772]*(-32)+in_buf[773]*(-38)+in_buf[774]*(-36)+in_buf[775]*(-39)+in_buf[776]*(-19)+in_buf[777]*(-32)+in_buf[778]*(-29)+in_buf[779]*(-22)+in_buf[780]*(3)+in_buf[781]*(0)+in_buf[782]*(-1)+in_buf[783]*(4);
assign in_buf_weight061=in_buf[0]*(4)+in_buf[1]*(1)+in_buf[2]*(0)+in_buf[3]*(4)+in_buf[4]*(4)+in_buf[5]*(2)+in_buf[6]*(1)+in_buf[7]*(4)+in_buf[8]*(-2)+in_buf[9]*(3)+in_buf[10]*(2)+in_buf[11]*(-1)+in_buf[12]*(-7)+in_buf[13]*(-8)+in_buf[14]*(15)+in_buf[15]*(5)+in_buf[16]*(0)+in_buf[17]*(3)+in_buf[18]*(3)+in_buf[19]*(3)+in_buf[20]*(-1)+in_buf[21]*(1)+in_buf[22]*(2)+in_buf[23]*(0)+in_buf[24]*(-1)+in_buf[25]*(-3)+in_buf[26]*(4)+in_buf[27]*(0)+in_buf[28]*(3)+in_buf[29]*(-3)+in_buf[30]*(2)+in_buf[31]*(4)+in_buf[32]*(-6)+in_buf[33]*(-9)+in_buf[34]*(-10)+in_buf[35]*(-8)+in_buf[36]*(-20)+in_buf[37]*(-8)+in_buf[38]*(-23)+in_buf[39]*(-31)+in_buf[40]*(-38)+in_buf[41]*(-39)+in_buf[42]*(-5)+in_buf[43]*(-18)+in_buf[44]*(-19)+in_buf[45]*(-27)+in_buf[46]*(-10)+in_buf[47]*(-25)+in_buf[48]*(-33)+in_buf[49]*(-14)+in_buf[50]*(3)+in_buf[51]*(0)+in_buf[52]*(0)+in_buf[53]*(1)+in_buf[54]*(-3)+in_buf[55]*(2)+in_buf[56]*(3)+in_buf[57]*(-2)+in_buf[58]*(-11)+in_buf[59]*(-8)+in_buf[60]*(-21)+in_buf[61]*(-18)+in_buf[62]*(-20)+in_buf[63]*(-25)+in_buf[64]*(-13)+in_buf[65]*(10)+in_buf[66]*(20)+in_buf[67]*(11)+in_buf[68]*(25)+in_buf[69]*(24)+in_buf[70]*(17)+in_buf[71]*(6)+in_buf[72]*(-6)+in_buf[73]*(-45)+in_buf[74]*(-47)+in_buf[75]*(-46)+in_buf[76]*(-55)+in_buf[77]*(-57)+in_buf[78]*(-47)+in_buf[79]*(-13)+in_buf[80]*(0)+in_buf[81]*(0)+in_buf[82]*(1)+in_buf[83]*(-2)+in_buf[84]*(0)+in_buf[85]*(0)+in_buf[86]*(17)+in_buf[87]*(2)+in_buf[88]*(-5)+in_buf[89]*(11)+in_buf[90]*(9)+in_buf[91]*(15)+in_buf[92]*(23)+in_buf[93]*(13)+in_buf[94]*(24)+in_buf[95]*(40)+in_buf[96]*(44)+in_buf[97]*(34)+in_buf[98]*(11)+in_buf[99]*(10)+in_buf[100]*(23)+in_buf[101]*(-19)+in_buf[102]*(-64)+in_buf[103]*(-55)+in_buf[104]*(-60)+in_buf[105]*(-81)+in_buf[106]*(-54)+in_buf[107]*(-48)+in_buf[108]*(-15)+in_buf[109]*(0)+in_buf[110]*(0)+in_buf[111]*(0)+in_buf[112]*(-2)+in_buf[113]*(5)+in_buf[114]*(8)+in_buf[115]*(30)+in_buf[116]*(42)+in_buf[117]*(34)+in_buf[118]*(17)+in_buf[119]*(13)+in_buf[120]*(38)+in_buf[121]*(27)+in_buf[122]*(19)+in_buf[123]*(20)+in_buf[124]*(24)+in_buf[125]*(19)+in_buf[126]*(11)+in_buf[127]*(14)+in_buf[128]*(2)+in_buf[129]*(-10)+in_buf[130]*(-14)+in_buf[131]*(-29)+in_buf[132]*(-43)+in_buf[133]*(-34)+in_buf[134]*(-22)+in_buf[135]*(-67)+in_buf[136]*(-28)+in_buf[137]*(0)+in_buf[138]*(-1)+in_buf[139]*(-1)+in_buf[140]*(0)+in_buf[141]*(2)+in_buf[142]*(-27)+in_buf[143]*(28)+in_buf[144]*(30)+in_buf[145]*(44)+in_buf[146]*(35)+in_buf[147]*(31)+in_buf[148]*(17)+in_buf[149]*(14)+in_buf[150]*(7)+in_buf[151]*(10)+in_buf[152]*(22)+in_buf[153]*(24)+in_buf[154]*(18)+in_buf[155]*(19)+in_buf[156]*(8)+in_buf[157]*(-5)+in_buf[158]*(-8)+in_buf[159]*(-25)+in_buf[160]*(-52)+in_buf[161]*(-51)+in_buf[162]*(-34)+in_buf[163]*(-81)+in_buf[164]*(-42)+in_buf[165]*(-5)+in_buf[166]*(-10)+in_buf[167]*(-3)+in_buf[168]*(-1)+in_buf[169]*(11)+in_buf[170]*(11)+in_buf[171]*(18)+in_buf[172]*(19)+in_buf[173]*(19)+in_buf[174]*(38)+in_buf[175]*(9)+in_buf[176]*(3)+in_buf[177]*(11)+in_buf[178]*(2)+in_buf[179]*(14)+in_buf[180]*(6)+in_buf[181]*(12)+in_buf[182]*(11)+in_buf[183]*(-4)+in_buf[184]*(11)+in_buf[185]*(5)+in_buf[186]*(0)+in_buf[187]*(-19)+in_buf[188]*(-22)+in_buf[189]*(-35)+in_buf[190]*(-56)+in_buf[191]*(-70)+in_buf[192]*(-42)+in_buf[193]*(-29)+in_buf[194]*(-25)+in_buf[195]*(6)+in_buf[196]*(5)+in_buf[197]*(34)+in_buf[198]*(3)+in_buf[199]*(31)+in_buf[200]*(48)+in_buf[201]*(14)+in_buf[202]*(18)+in_buf[203]*(10)+in_buf[204]*(-9)+in_buf[205]*(5)+in_buf[206]*(2)+in_buf[207]*(-4)+in_buf[208]*(0)+in_buf[209]*(5)+in_buf[210]*(6)+in_buf[211]*(0)+in_buf[212]*(8)+in_buf[213]*(27)+in_buf[214]*(1)+in_buf[215]*(-17)+in_buf[216]*(-27)+in_buf[217]*(-65)+in_buf[218]*(-91)+in_buf[219]*(-81)+in_buf[220]*(-42)+in_buf[221]*(-29)+in_buf[222]*(-15)+in_buf[223]*(-3)+in_buf[224]*(-11)+in_buf[225]*(4)+in_buf[226]*(28)+in_buf[227]*(29)+in_buf[228]*(33)+in_buf[229]*(13)+in_buf[230]*(-6)+in_buf[231]*(1)+in_buf[232]*(-20)+in_buf[233]*(-18)+in_buf[234]*(-11)+in_buf[235]*(-31)+in_buf[236]*(-21)+in_buf[237]*(0)+in_buf[238]*(17)+in_buf[239]*(35)+in_buf[240]*(27)+in_buf[241]*(31)+in_buf[242]*(1)+in_buf[243]*(-15)+in_buf[244]*(-41)+in_buf[245]*(-75)+in_buf[246]*(-73)+in_buf[247]*(-69)+in_buf[248]*(-52)+in_buf[249]*(-38)+in_buf[250]*(-6)+in_buf[251]*(0)+in_buf[252]*(16)+in_buf[253]*(15)+in_buf[254]*(28)+in_buf[255]*(10)+in_buf[256]*(38)+in_buf[257]*(22)+in_buf[258]*(-6)+in_buf[259]*(-6)+in_buf[260]*(-30)+in_buf[261]*(-30)+in_buf[262]*(-47)+in_buf[263]*(-37)+in_buf[264]*(-16)+in_buf[265]*(0)+in_buf[266]*(31)+in_buf[267]*(55)+in_buf[268]*(52)+in_buf[269]*(19)+in_buf[270]*(-4)+in_buf[271]*(-26)+in_buf[272]*(-59)+in_buf[273]*(-76)+in_buf[274]*(-64)+in_buf[275]*(-59)+in_buf[276]*(-62)+in_buf[277]*(-37)+in_buf[278]*(-23)+in_buf[279]*(-14)+in_buf[280]*(15)+in_buf[281]*(7)+in_buf[282]*(24)+in_buf[283]*(2)+in_buf[284]*(1)+in_buf[285]*(-5)+in_buf[286]*(-18)+in_buf[287]*(-32)+in_buf[288]*(-55)+in_buf[289]*(-56)+in_buf[290]*(-33)+in_buf[291]*(-19)+in_buf[292]*(-8)+in_buf[293]*(23)+in_buf[294]*(31)+in_buf[295]*(32)+in_buf[296]*(32)+in_buf[297]*(21)+in_buf[298]*(-15)+in_buf[299]*(-39)+in_buf[300]*(-64)+in_buf[301]*(-43)+in_buf[302]*(-25)+in_buf[303]*(-21)+in_buf[304]*(-36)+in_buf[305]*(24)+in_buf[306]*(25)+in_buf[307]*(25)+in_buf[308]*(7)+in_buf[309]*(32)+in_buf[310]*(-5)+in_buf[311]*(5)+in_buf[312]*(-2)+in_buf[313]*(-29)+in_buf[314]*(-38)+in_buf[315]*(-37)+in_buf[316]*(-39)+in_buf[317]*(-19)+in_buf[318]*(3)+in_buf[319]*(9)+in_buf[320]*(14)+in_buf[321]*(24)+in_buf[322]*(32)+in_buf[323]*(19)+in_buf[324]*(4)+in_buf[325]*(-5)+in_buf[326]*(-22)+in_buf[327]*(-33)+in_buf[328]*(-37)+in_buf[329]*(-47)+in_buf[330]*(-14)+in_buf[331]*(4)+in_buf[332]*(-9)+in_buf[333]*(19)+in_buf[334]*(15)+in_buf[335]*(32)+in_buf[336]*(6)+in_buf[337]*(20)+in_buf[338]*(13)+in_buf[339]*(-6)+in_buf[340]*(-38)+in_buf[341]*(-31)+in_buf[342]*(-33)+in_buf[343]*(-22)+in_buf[344]*(-6)+in_buf[345]*(19)+in_buf[346]*(27)+in_buf[347]*(18)+in_buf[348]*(24)+in_buf[349]*(14)+in_buf[350]*(18)+in_buf[351]*(7)+in_buf[352]*(0)+in_buf[353]*(-18)+in_buf[354]*(-28)+in_buf[355]*(-36)+in_buf[356]*(-23)+in_buf[357]*(-24)+in_buf[358]*(-25)+in_buf[359]*(-6)+in_buf[360]*(30)+in_buf[361]*(34)+in_buf[362]*(-4)+in_buf[363]*(30)+in_buf[364]*(-6)+in_buf[365]*(1)+in_buf[366]*(23)+in_buf[367]*(-10)+in_buf[368]*(-47)+in_buf[369]*(-56)+in_buf[370]*(-1)+in_buf[371]*(3)+in_buf[372]*(20)+in_buf[373]*(30)+in_buf[374]*(22)+in_buf[375]*(10)+in_buf[376]*(5)+in_buf[377]*(11)+in_buf[378]*(11)+in_buf[379]*(-2)+in_buf[380]*(6)+in_buf[381]*(-7)+in_buf[382]*(-11)+in_buf[383]*(-29)+in_buf[384]*(-6)+in_buf[385]*(10)+in_buf[386]*(-7)+in_buf[387]*(-7)+in_buf[388]*(20)+in_buf[389]*(43)+in_buf[390]*(6)+in_buf[391]*(7)+in_buf[392]*(-13)+in_buf[393]*(7)+in_buf[394]*(19)+in_buf[395]*(17)+in_buf[396]*(-13)+in_buf[397]*(-29)+in_buf[398]*(-18)+in_buf[399]*(6)+in_buf[400]*(24)+in_buf[401]*(12)+in_buf[402]*(-2)+in_buf[403]*(-7)+in_buf[404]*(-5)+in_buf[405]*(-2)+in_buf[406]*(8)+in_buf[407]*(7)+in_buf[408]*(10)+in_buf[409]*(6)+in_buf[410]*(-3)+in_buf[411]*(3)+in_buf[412]*(5)+in_buf[413]*(38)+in_buf[414]*(15)+in_buf[415]*(20)+in_buf[416]*(25)+in_buf[417]*(37)+in_buf[418]*(15)+in_buf[419]*(-3)+in_buf[420]*(-11)+in_buf[421]*(7)+in_buf[422]*(16)+in_buf[423]*(22)+in_buf[424]*(0)+in_buf[425]*(-25)+in_buf[426]*(-11)+in_buf[427]*(16)+in_buf[428]*(23)+in_buf[429]*(3)+in_buf[430]*(-21)+in_buf[431]*(-14)+in_buf[432]*(-13)+in_buf[433]*(0)+in_buf[434]*(11)+in_buf[435]*(6)+in_buf[436]*(13)+in_buf[437]*(3)+in_buf[438]*(-14)+in_buf[439]*(3)+in_buf[440]*(25)+in_buf[441]*(35)+in_buf[442]*(34)+in_buf[443]*(31)+in_buf[444]*(52)+in_buf[445]*(5)+in_buf[446]*(58)+in_buf[447]*(25)+in_buf[448]*(0)+in_buf[449]*(3)+in_buf[450]*(12)+in_buf[451]*(8)+in_buf[452]*(0)+in_buf[453]*(-27)+in_buf[454]*(8)+in_buf[455]*(34)+in_buf[456]*(28)+in_buf[457]*(21)+in_buf[458]*(-23)+in_buf[459]*(-18)+in_buf[460]*(-9)+in_buf[461]*(-2)+in_buf[462]*(7)+in_buf[463]*(-5)+in_buf[464]*(9)+in_buf[465]*(-2)+in_buf[466]*(-2)+in_buf[467]*(11)+in_buf[468]*(16)+in_buf[469]*(26)+in_buf[470]*(13)+in_buf[471]*(32)+in_buf[472]*(56)+in_buf[473]*(-18)+in_buf[474]*(25)+in_buf[475]*(25)+in_buf[476]*(1)+in_buf[477]*(7)+in_buf[478]*(21)+in_buf[479]*(3)+in_buf[480]*(1)+in_buf[481]*(-21)+in_buf[482]*(-9)+in_buf[483]*(19)+in_buf[484]*(11)+in_buf[485]*(-7)+in_buf[486]*(-29)+in_buf[487]*(-17)+in_buf[488]*(-2)+in_buf[489]*(24)+in_buf[490]*(10)+in_buf[491]*(-8)+in_buf[492]*(1)+in_buf[493]*(-1)+in_buf[494]*(-7)+in_buf[495]*(4)+in_buf[496]*(5)+in_buf[497]*(23)+in_buf[498]*(22)+in_buf[499]*(38)+in_buf[500]*(41)+in_buf[501]*(2)+in_buf[502]*(22)+in_buf[503]*(-22)+in_buf[504]*(-44)+in_buf[505]*(17)+in_buf[506]*(32)+in_buf[507]*(0)+in_buf[508]*(9)+in_buf[509]*(12)+in_buf[510]*(-3)+in_buf[511]*(-9)+in_buf[512]*(2)+in_buf[513]*(-9)+in_buf[514]*(-22)+in_buf[515]*(-21)+in_buf[516]*(-12)+in_buf[517]*(15)+in_buf[518]*(-4)+in_buf[519]*(-16)+in_buf[520]*(5)+in_buf[521]*(0)+in_buf[522]*(0)+in_buf[523]*(7)+in_buf[524]*(10)+in_buf[525]*(24)+in_buf[526]*(26)+in_buf[527]*(24)+in_buf[528]*(17)+in_buf[529]*(-9)+in_buf[530]*(30)+in_buf[531]*(12)+in_buf[532]*(25)+in_buf[533]*(-32)+in_buf[534]*(-2)+in_buf[535]*(9)+in_buf[536]*(4)+in_buf[537]*(10)+in_buf[538]*(-12)+in_buf[539]*(-11)+in_buf[540]*(-10)+in_buf[541]*(-11)+in_buf[542]*(-20)+in_buf[543]*(-31)+in_buf[544]*(-9)+in_buf[545]*(5)+in_buf[546]*(2)+in_buf[547]*(-3)+in_buf[548]*(7)+in_buf[549]*(3)+in_buf[550]*(0)+in_buf[551]*(-1)+in_buf[552]*(-1)+in_buf[553]*(19)+in_buf[554]*(10)+in_buf[555]*(2)+in_buf[556]*(-12)+in_buf[557]*(0)+in_buf[558]*(12)+in_buf[559]*(5)+in_buf[560]*(-2)+in_buf[561]*(-25)+in_buf[562]*(0)+in_buf[563]*(5)+in_buf[564]*(-27)+in_buf[565]*(-3)+in_buf[566]*(6)+in_buf[567]*(-2)+in_buf[568]*(-2)+in_buf[569]*(9)+in_buf[570]*(-5)+in_buf[571]*(-12)+in_buf[572]*(-3)+in_buf[573]*(-6)+in_buf[574]*(11)+in_buf[575]*(-9)+in_buf[576]*(3)+in_buf[577]*(-4)+in_buf[578]*(3)+in_buf[579]*(-6)+in_buf[580]*(1)+in_buf[581]*(-2)+in_buf[582]*(-7)+in_buf[583]*(4)+in_buf[584]*(3)+in_buf[585]*(-14)+in_buf[586]*(9)+in_buf[587]*(13)+in_buf[588]*(29)+in_buf[589]*(16)+in_buf[590]*(42)+in_buf[591]*(10)+in_buf[592]*(-29)+in_buf[593]*(-12)+in_buf[594]*(7)+in_buf[595]*(-7)+in_buf[596]*(-6)+in_buf[597]*(-9)+in_buf[598]*(5)+in_buf[599]*(-2)+in_buf[600]*(-3)+in_buf[601]*(-8)+in_buf[602]*(-5)+in_buf[603]*(2)+in_buf[604]*(1)+in_buf[605]*(-4)+in_buf[606]*(-5)+in_buf[607]*(-5)+in_buf[608]*(-13)+in_buf[609]*(-25)+in_buf[610]*(-4)+in_buf[611]*(-10)+in_buf[612]*(-22)+in_buf[613]*(0)+in_buf[614]*(-30)+in_buf[615]*(-2)+in_buf[616]*(21)+in_buf[617]*(38)+in_buf[618]*(25)+in_buf[619]*(20)+in_buf[620]*(27)+in_buf[621]*(18)+in_buf[622]*(14)+in_buf[623]*(-1)+in_buf[624]*(-7)+in_buf[625]*(-10)+in_buf[626]*(1)+in_buf[627]*(-5)+in_buf[628]*(-8)+in_buf[629]*(0)+in_buf[630]*(1)+in_buf[631]*(-1)+in_buf[632]*(-8)+in_buf[633]*(-5)+in_buf[634]*(8)+in_buf[635]*(8)+in_buf[636]*(5)+in_buf[637]*(-1)+in_buf[638]*(1)+in_buf[639]*(-25)+in_buf[640]*(-27)+in_buf[641]*(-10)+in_buf[642]*(-2)+in_buf[643]*(-3)+in_buf[644]*(0)+in_buf[645]*(-1)+in_buf[646]*(16)+in_buf[647]*(13)+in_buf[648]*(36)+in_buf[649]*(27)+in_buf[650]*(11)+in_buf[651]*(20)+in_buf[652]*(5)+in_buf[653]*(3)+in_buf[654]*(12)+in_buf[655]*(13)+in_buf[656]*(6)+in_buf[657]*(9)+in_buf[658]*(-10)+in_buf[659]*(-4)+in_buf[660]*(-8)+in_buf[661]*(0)+in_buf[662]*(12)+in_buf[663]*(15)+in_buf[664]*(18)+in_buf[665]*(-5)+in_buf[666]*(-17)+in_buf[667]*(-41)+in_buf[668]*(-20)+in_buf[669]*(-13)+in_buf[670]*(10)+in_buf[671]*(4)+in_buf[672]*(3)+in_buf[673]*(1)+in_buf[674]*(20)+in_buf[675]*(7)+in_buf[676]*(26)+in_buf[677]*(26)+in_buf[678]*(25)+in_buf[679]*(26)+in_buf[680]*(15)+in_buf[681]*(13)+in_buf[682]*(10)+in_buf[683]*(14)+in_buf[684]*(0)+in_buf[685]*(2)+in_buf[686]*(11)+in_buf[687]*(-12)+in_buf[688]*(-11)+in_buf[689]*(2)+in_buf[690]*(7)+in_buf[691]*(13)+in_buf[692]*(3)+in_buf[693]*(26)+in_buf[694]*(4)+in_buf[695]*(3)+in_buf[696]*(0)+in_buf[697]*(2)+in_buf[698]*(26)+in_buf[699]*(-3)+in_buf[700]*(0)+in_buf[701]*(0)+in_buf[702]*(8)+in_buf[703]*(-8)+in_buf[704]*(21)+in_buf[705]*(39)+in_buf[706]*(64)+in_buf[707]*(62)+in_buf[708]*(62)+in_buf[709]*(20)+in_buf[710]*(12)+in_buf[711]*(16)+in_buf[712]*(7)+in_buf[713]*(3)+in_buf[714]*(0)+in_buf[715]*(-27)+in_buf[716]*(-34)+in_buf[717]*(-22)+in_buf[718]*(2)+in_buf[719]*(0)+in_buf[720]*(25)+in_buf[721]*(-2)+in_buf[722]*(16)+in_buf[723]*(1)+in_buf[724]*(-13)+in_buf[725]*(-3)+in_buf[726]*(4)+in_buf[727]*(2)+in_buf[728]*(-3)+in_buf[729]*(1)+in_buf[730]*(-2)+in_buf[731]*(-2)+in_buf[732]*(6)+in_buf[733]*(-8)+in_buf[734]*(-30)+in_buf[735]*(-27)+in_buf[736]*(-30)+in_buf[737]*(-31)+in_buf[738]*(0)+in_buf[739]*(25)+in_buf[740]*(1)+in_buf[741]*(-1)+in_buf[742]*(-5)+in_buf[743]*(1)+in_buf[744]*(0)+in_buf[745]*(16)+in_buf[746]*(23)+in_buf[747]*(11)+in_buf[748]*(8)+in_buf[749]*(-32)+in_buf[750]*(-28)+in_buf[751]*(-18)+in_buf[752]*(1)+in_buf[753]*(-2)+in_buf[754]*(-3)+in_buf[755]*(-1)+in_buf[756]*(2)+in_buf[757]*(-3)+in_buf[758]*(-3)+in_buf[759]*(0)+in_buf[760]*(5)+in_buf[761]*(0)+in_buf[762]*(-10)+in_buf[763]*(-5)+in_buf[764]*(-5)+in_buf[765]*(-6)+in_buf[766]*(-36)+in_buf[767]*(-23)+in_buf[768]*(-14)+in_buf[769]*(-16)+in_buf[770]*(-52)+in_buf[771]*(-22)+in_buf[772]*(-4)+in_buf[773]*(-8)+in_buf[774]*(-4)+in_buf[775]*(7)+in_buf[776]*(3)+in_buf[777]*(-2)+in_buf[778]*(2)+in_buf[779]*(0)+in_buf[780]*(-2)+in_buf[781]*(-2)+in_buf[782]*(1)+in_buf[783]*(4);
assign in_buf_weight062=in_buf[0]*(0)+in_buf[1]*(1)+in_buf[2]*(0)+in_buf[3]*(3)+in_buf[4]*(-1)+in_buf[5]*(-2)+in_buf[6]*(-3)+in_buf[7]*(2)+in_buf[8]*(-2)+in_buf[9]*(2)+in_buf[10]*(1)+in_buf[11]*(0)+in_buf[12]*(4)+in_buf[13]*(6)+in_buf[14]*(0)+in_buf[15]*(0)+in_buf[16]*(-3)+in_buf[17]*(-1)+in_buf[18]*(4)+in_buf[19]*(-1)+in_buf[20]*(-2)+in_buf[21]*(-2)+in_buf[22]*(0)+in_buf[23]*(-2)+in_buf[24]*(3)+in_buf[25]*(0)+in_buf[26]*(-1)+in_buf[27]*(-3)+in_buf[28]*(-3)+in_buf[29]*(0)+in_buf[30]*(0)+in_buf[31]*(-3)+in_buf[32]*(4)+in_buf[33]*(5)+in_buf[34]*(3)+in_buf[35]*(2)+in_buf[36]*(6)+in_buf[37]*(6)+in_buf[38]*(5)+in_buf[39]*(12)+in_buf[40]*(5)+in_buf[41]*(9)+in_buf[42]*(1)+in_buf[43]*(1)+in_buf[44]*(3)+in_buf[45]*(0)+in_buf[46]*(-1)+in_buf[47]*(1)+in_buf[48]*(0)+in_buf[49]*(0)+in_buf[50]*(-1)+in_buf[51]*(5)+in_buf[52]*(4)+in_buf[53]*(1)+in_buf[54]*(-2)+in_buf[55]*(1)+in_buf[56]*(-2)+in_buf[57]*(-3)+in_buf[58]*(-1)+in_buf[59]*(3)+in_buf[60]*(-8)+in_buf[61]*(3)+in_buf[62]*(0)+in_buf[63]*(11)+in_buf[64]*(0)+in_buf[65]*(-11)+in_buf[66]*(-15)+in_buf[67]*(1)+in_buf[68]*(30)+in_buf[69]*(20)+in_buf[70]*(-17)+in_buf[71]*(-39)+in_buf[72]*(-37)+in_buf[73]*(2)+in_buf[74]*(7)+in_buf[75]*(-34)+in_buf[76]*(-38)+in_buf[77]*(-10)+in_buf[78]*(-15)+in_buf[79]*(-1)+in_buf[80]*(-8)+in_buf[81]*(-1)+in_buf[82]*(0)+in_buf[83]*(0)+in_buf[84]*(0)+in_buf[85]*(2)+in_buf[86]*(-23)+in_buf[87]*(0)+in_buf[88]*(-2)+in_buf[89]*(-4)+in_buf[90]*(-5)+in_buf[91]*(-4)+in_buf[92]*(-11)+in_buf[93]*(-5)+in_buf[94]*(-12)+in_buf[95]*(-1)+in_buf[96]*(34)+in_buf[97]*(30)+in_buf[98]*(-3)+in_buf[99]*(-30)+in_buf[100]*(-34)+in_buf[101]*(-17)+in_buf[102]*(11)+in_buf[103]*(-34)+in_buf[104]*(-51)+in_buf[105]*(-35)+in_buf[106]*(-16)+in_buf[107]*(8)+in_buf[108]*(1)+in_buf[109]*(-22)+in_buf[110]*(-24)+in_buf[111]*(0)+in_buf[112]*(-3)+in_buf[113]*(4)+in_buf[114]*(-16)+in_buf[115]*(-2)+in_buf[116]*(11)+in_buf[117]*(-12)+in_buf[118]*(-11)+in_buf[119]*(-1)+in_buf[120]*(3)+in_buf[121]*(14)+in_buf[122]*(4)+in_buf[123]*(29)+in_buf[124]*(31)+in_buf[125]*(11)+in_buf[126]*(-7)+in_buf[127]*(3)+in_buf[128]*(12)+in_buf[129]*(1)+in_buf[130]*(3)+in_buf[131]*(-7)+in_buf[132]*(-19)+in_buf[133]*(-11)+in_buf[134]*(-8)+in_buf[135]*(-23)+in_buf[136]*(-24)+in_buf[137]*(-7)+in_buf[138]*(20)+in_buf[139]*(14)+in_buf[140]*(0)+in_buf[141]*(1)+in_buf[142]*(18)+in_buf[143]*(44)+in_buf[144]*(32)+in_buf[145]*(-8)+in_buf[146]*(-12)+in_buf[147]*(-3)+in_buf[148]*(-10)+in_buf[149]*(-8)+in_buf[150]*(11)+in_buf[151]*(14)+in_buf[152]*(9)+in_buf[153]*(9)+in_buf[154]*(10)+in_buf[155]*(7)+in_buf[156]*(15)+in_buf[157]*(12)+in_buf[158]*(3)+in_buf[159]*(6)+in_buf[160]*(21)+in_buf[161]*(23)+in_buf[162]*(23)+in_buf[163]*(-6)+in_buf[164]*(-5)+in_buf[165]*(14)+in_buf[166]*(36)+in_buf[167]*(3)+in_buf[168]*(-2)+in_buf[169]*(5)+in_buf[170]*(4)+in_buf[171]*(16)+in_buf[172]*(-10)+in_buf[173]*(-14)+in_buf[174]*(-14)+in_buf[175]*(-3)+in_buf[176]*(0)+in_buf[177]*(-2)+in_buf[178]*(12)+in_buf[179]*(10)+in_buf[180]*(6)+in_buf[181]*(-2)+in_buf[182]*(-1)+in_buf[183]*(4)+in_buf[184]*(-3)+in_buf[185]*(-2)+in_buf[186]*(5)+in_buf[187]*(-6)+in_buf[188]*(-12)+in_buf[189]*(2)+in_buf[190]*(14)+in_buf[191]*(8)+in_buf[192]*(13)+in_buf[193]*(-7)+in_buf[194]*(41)+in_buf[195]*(32)+in_buf[196]*(-16)+in_buf[197]*(-3)+in_buf[198]*(0)+in_buf[199]*(-10)+in_buf[200]*(20)+in_buf[201]*(19)+in_buf[202]*(-4)+in_buf[203]*(-1)+in_buf[204]*(7)+in_buf[205]*(5)+in_buf[206]*(11)+in_buf[207]*(6)+in_buf[208]*(-3)+in_buf[209]*(-1)+in_buf[210]*(-1)+in_buf[211]*(0)+in_buf[212]*(5)+in_buf[213]*(-12)+in_buf[214]*(12)+in_buf[215]*(3)+in_buf[216]*(-11)+in_buf[217]*(4)+in_buf[218]*(19)+in_buf[219]*(3)+in_buf[220]*(-14)+in_buf[221]*(-24)+in_buf[222]*(-1)+in_buf[223]*(24)+in_buf[224]*(-14)+in_buf[225]*(-29)+in_buf[226]*(-12)+in_buf[227]*(18)+in_buf[228]*(33)+in_buf[229]*(5)+in_buf[230]*(-1)+in_buf[231]*(0)+in_buf[232]*(-9)+in_buf[233]*(-4)+in_buf[234]*(6)+in_buf[235]*(3)+in_buf[236]*(5)+in_buf[237]*(2)+in_buf[238]*(-3)+in_buf[239]*(-11)+in_buf[240]*(10)+in_buf[241]*(12)+in_buf[242]*(5)+in_buf[243]*(15)+in_buf[244]*(7)+in_buf[245]*(-10)+in_buf[246]*(15)+in_buf[247]*(4)+in_buf[248]*(-21)+in_buf[249]*(-14)+in_buf[250]*(9)+in_buf[251]*(18)+in_buf[252]*(-16)+in_buf[253]*(-13)+in_buf[254]*(5)+in_buf[255]*(24)+in_buf[256]*(16)+in_buf[257]*(-5)+in_buf[258]*(-7)+in_buf[259]*(5)+in_buf[260]*(10)+in_buf[261]*(2)+in_buf[262]*(7)+in_buf[263]*(-2)+in_buf[264]*(-1)+in_buf[265]*(6)+in_buf[266]*(0)+in_buf[267]*(-2)+in_buf[268]*(17)+in_buf[269]*(6)+in_buf[270]*(5)+in_buf[271]*(15)+in_buf[272]*(0)+in_buf[273]*(-10)+in_buf[274]*(6)+in_buf[275]*(26)+in_buf[276]*(16)+in_buf[277]*(33)+in_buf[278]*(1)+in_buf[279]*(-24)+in_buf[280]*(-15)+in_buf[281]*(2)+in_buf[282]*(5)+in_buf[283]*(13)+in_buf[284]*(6)+in_buf[285]*(-1)+in_buf[286]*(1)+in_buf[287]*(0)+in_buf[288]*(13)+in_buf[289]*(0)+in_buf[290]*(10)+in_buf[291]*(-1)+in_buf[292]*(-2)+in_buf[293]*(15)+in_buf[294]*(17)+in_buf[295]*(9)+in_buf[296]*(4)+in_buf[297]*(4)+in_buf[298]*(12)+in_buf[299]*(20)+in_buf[300]*(16)+in_buf[301]*(3)+in_buf[302]*(4)+in_buf[303]*(31)+in_buf[304]*(28)+in_buf[305]*(-5)+in_buf[306]*(2)+in_buf[307]*(-19)+in_buf[308]*(-27)+in_buf[309]*(-13)+in_buf[310]*(-37)+in_buf[311]*(3)+in_buf[312]*(24)+in_buf[313]*(-6)+in_buf[314]*(1)+in_buf[315]*(4)+in_buf[316]*(-3)+in_buf[317]*(-2)+in_buf[318]*(-14)+in_buf[319]*(-13)+in_buf[320]*(-7)+in_buf[321]*(9)+in_buf[322]*(10)+in_buf[323]*(-8)+in_buf[324]*(-23)+in_buf[325]*(-14)+in_buf[326]*(0)+in_buf[327]*(6)+in_buf[328]*(0)+in_buf[329]*(18)+in_buf[330]*(0)+in_buf[331]*(-1)+in_buf[332]*(4)+in_buf[333]*(25)+in_buf[334]*(52)+in_buf[335]*(6)+in_buf[336]*(-19)+in_buf[337]*(-31)+in_buf[338]*(-45)+in_buf[339]*(8)+in_buf[340]*(-1)+in_buf[341]*(-21)+in_buf[342]*(-8)+in_buf[343]*(11)+in_buf[344]*(7)+in_buf[345]*(14)+in_buf[346]*(-14)+in_buf[347]*(-18)+in_buf[348]*(-8)+in_buf[349]*(-13)+in_buf[350]*(-16)+in_buf[351]*(-31)+in_buf[352]*(-33)+in_buf[353]*(-18)+in_buf[354]*(-14)+in_buf[355]*(0)+in_buf[356]*(8)+in_buf[357]*(12)+in_buf[358]*(-5)+in_buf[359]*(-19)+in_buf[360]*(27)+in_buf[361]*(60)+in_buf[362]*(43)+in_buf[363]*(10)+in_buf[364]*(27)+in_buf[365]*(-38)+in_buf[366]*(-49)+in_buf[367]*(14)+in_buf[368]*(-13)+in_buf[369]*(-22)+in_buf[370]*(1)+in_buf[371]*(0)+in_buf[372]*(-2)+in_buf[373]*(4)+in_buf[374]*(-26)+in_buf[375]*(-10)+in_buf[376]*(0)+in_buf[377]*(-6)+in_buf[378]*(-12)+in_buf[379]*(-28)+in_buf[380]*(-34)+in_buf[381]*(-16)+in_buf[382]*(-6)+in_buf[383]*(-4)+in_buf[384]*(-4)+in_buf[385]*(-10)+in_buf[386]*(-8)+in_buf[387]*(-17)+in_buf[388]*(1)+in_buf[389]*(34)+in_buf[390]*(29)+in_buf[391]*(11)+in_buf[392]*(14)+in_buf[393]*(-33)+in_buf[394]*(-37)+in_buf[395]*(-4)+in_buf[396]*(-31)+in_buf[397]*(-26)+in_buf[398]*(-7)+in_buf[399]*(-13)+in_buf[400]*(-12)+in_buf[401]*(-23)+in_buf[402]*(-29)+in_buf[403]*(-4)+in_buf[404]*(-2)+in_buf[405]*(0)+in_buf[406]*(-11)+in_buf[407]*(-30)+in_buf[408]*(-30)+in_buf[409]*(-13)+in_buf[410]*(-10)+in_buf[411]*(-33)+in_buf[412]*(-6)+in_buf[413]*(-3)+in_buf[414]*(-15)+in_buf[415]*(-37)+in_buf[416]*(-15)+in_buf[417]*(-4)+in_buf[418]*(27)+in_buf[419]*(21)+in_buf[420]*(12)+in_buf[421]*(-7)+in_buf[422]*(-25)+in_buf[423]*(-12)+in_buf[424]*(-34)+in_buf[425]*(-13)+in_buf[426]*(1)+in_buf[427]*(0)+in_buf[428]*(0)+in_buf[429]*(1)+in_buf[430]*(-13)+in_buf[431]*(5)+in_buf[432]*(13)+in_buf[433]*(14)+in_buf[434]*(9)+in_buf[435]*(-23)+in_buf[436]*(-15)+in_buf[437]*(-25)+in_buf[438]*(-28)+in_buf[439]*(-29)+in_buf[440]*(-9)+in_buf[441]*(-11)+in_buf[442]*(-37)+in_buf[443]*(-24)+in_buf[444]*(0)+in_buf[445]*(-29)+in_buf[446]*(-9)+in_buf[447]*(15)+in_buf[448]*(-13)+in_buf[449]*(1)+in_buf[450]*(2)+in_buf[451]*(5)+in_buf[452]*(-15)+in_buf[453]*(-18)+in_buf[454]*(-30)+in_buf[455]*(-15)+in_buf[456]*(-1)+in_buf[457]*(12)+in_buf[458]*(16)+in_buf[459]*(21)+in_buf[460]*(4)+in_buf[461]*(21)+in_buf[462]*(9)+in_buf[463]*(-15)+in_buf[464]*(-14)+in_buf[465]*(-29)+in_buf[466]*(-25)+in_buf[467]*(-17)+in_buf[468]*(-21)+in_buf[469]*(-14)+in_buf[470]*(-17)+in_buf[471]*(-4)+in_buf[472]*(-13)+in_buf[473]*(-3)+in_buf[474]*(19)+in_buf[475]*(26)+in_buf[476]*(3)+in_buf[477]*(-9)+in_buf[478]*(-6)+in_buf[479]*(6)+in_buf[480]*(0)+in_buf[481]*(-17)+in_buf[482]*(-26)+in_buf[483]*(-17)+in_buf[484]*(-9)+in_buf[485]*(-1)+in_buf[486]*(20)+in_buf[487]*(10)+in_buf[488]*(8)+in_buf[489]*(13)+in_buf[490]*(9)+in_buf[491]*(-16)+in_buf[492]*(-19)+in_buf[493]*(-24)+in_buf[494]*(-34)+in_buf[495]*(-4)+in_buf[496]*(-6)+in_buf[497]*(-8)+in_buf[498]*(3)+in_buf[499]*(-12)+in_buf[500]*(-11)+in_buf[501]*(-7)+in_buf[502]*(-5)+in_buf[503]*(35)+in_buf[504]*(0)+in_buf[505]*(7)+in_buf[506]*(-8)+in_buf[507]*(3)+in_buf[508]*(7)+in_buf[509]*(-6)+in_buf[510]*(-24)+in_buf[511]*(-11)+in_buf[512]*(-12)+in_buf[513]*(-3)+in_buf[514]*(-3)+in_buf[515]*(-11)+in_buf[516]*(1)+in_buf[517]*(-1)+in_buf[518]*(-14)+in_buf[519]*(-12)+in_buf[520]*(-7)+in_buf[521]*(-25)+in_buf[522]*(-28)+in_buf[523]*(-10)+in_buf[524]*(-8)+in_buf[525]*(-4)+in_buf[526]*(2)+in_buf[527]*(9)+in_buf[528]*(-1)+in_buf[529]*(0)+in_buf[530]*(-9)+in_buf[531]*(32)+in_buf[532]*(17)+in_buf[533]*(3)+in_buf[534]*(24)+in_buf[535]*(6)+in_buf[536]*(3)+in_buf[537]*(-6)+in_buf[538]*(-14)+in_buf[539]*(-2)+in_buf[540]*(-7)+in_buf[541]*(-12)+in_buf[542]*(0)+in_buf[543]*(-15)+in_buf[544]*(-1)+in_buf[545]*(2)+in_buf[546]*(-11)+in_buf[547]*(0)+in_buf[548]*(3)+in_buf[549]*(0)+in_buf[550]*(3)+in_buf[551]*(-4)+in_buf[552]*(4)+in_buf[553]*(7)+in_buf[554]*(27)+in_buf[555]*(58)+in_buf[556]*(0)+in_buf[557]*(24)+in_buf[558]*(52)+in_buf[559]*(26)+in_buf[560]*(0)+in_buf[561]*(5)+in_buf[562]*(38)+in_buf[563]*(35)+in_buf[564]*(22)+in_buf[565]*(-4)+in_buf[566]*(17)+in_buf[567]*(15)+in_buf[568]*(9)+in_buf[569]*(4)+in_buf[570]*(-9)+in_buf[571]*(0)+in_buf[572]*(8)+in_buf[573]*(7)+in_buf[574]*(7)+in_buf[575]*(20)+in_buf[576]*(14)+in_buf[577]*(22)+in_buf[578]*(28)+in_buf[579]*(24)+in_buf[580]*(37)+in_buf[581]*(45)+in_buf[582]*(50)+in_buf[583]*(60)+in_buf[584]*(-2)+in_buf[585]*(44)+in_buf[586]*(36)+in_buf[587]*(14)+in_buf[588]*(3)+in_buf[589]*(14)+in_buf[590]*(39)+in_buf[591]*(57)+in_buf[592]*(25)+in_buf[593]*(8)+in_buf[594]*(27)+in_buf[595]*(24)+in_buf[596]*(4)+in_buf[597]*(16)+in_buf[598]*(-2)+in_buf[599]*(13)+in_buf[600]*(6)+in_buf[601]*(27)+in_buf[602]*(43)+in_buf[603]*(49)+in_buf[604]*(30)+in_buf[605]*(44)+in_buf[606]*(41)+in_buf[607]*(43)+in_buf[608]*(41)+in_buf[609]*(17)+in_buf[610]*(41)+in_buf[611]*(50)+in_buf[612]*(25)+in_buf[613]*(49)+in_buf[614]*(37)+in_buf[615]*(-2)+in_buf[616]*(2)+in_buf[617]*(-9)+in_buf[618]*(48)+in_buf[619]*(58)+in_buf[620]*(19)+in_buf[621]*(30)+in_buf[622]*(35)+in_buf[623]*(23)+in_buf[624]*(31)+in_buf[625]*(35)+in_buf[626]*(10)+in_buf[627]*(32)+in_buf[628]*(26)+in_buf[629]*(35)+in_buf[630]*(33)+in_buf[631]*(28)+in_buf[632]*(33)+in_buf[633]*(45)+in_buf[634]*(27)+in_buf[635]*(34)+in_buf[636]*(29)+in_buf[637]*(11)+in_buf[638]*(20)+in_buf[639]*(43)+in_buf[640]*(52)+in_buf[641]*(20)+in_buf[642]*(3)+in_buf[643]*(-2)+in_buf[644]*(0)+in_buf[645]*(-3)+in_buf[646]*(31)+in_buf[647]*(40)+in_buf[648]*(18)+in_buf[649]*(15)+in_buf[650]*(29)+in_buf[651]*(21)+in_buf[652]*(42)+in_buf[653]*(44)+in_buf[654]*(33)+in_buf[655]*(41)+in_buf[656]*(41)+in_buf[657]*(35)+in_buf[658]*(25)+in_buf[659]*(35)+in_buf[660]*(42)+in_buf[661]*(39)+in_buf[662]*(27)+in_buf[663]*(31)+in_buf[664]*(31)+in_buf[665]*(19)+in_buf[666]*(50)+in_buf[667]*(47)+in_buf[668]*(43)+in_buf[669]*(27)+in_buf[670]*(9)+in_buf[671]*(5)+in_buf[672]*(4)+in_buf[673]*(3)+in_buf[674]*(-7)+in_buf[675]*(8)+in_buf[676]*(0)+in_buf[677]*(1)+in_buf[678]*(8)+in_buf[679]*(6)+in_buf[680]*(11)+in_buf[681]*(28)+in_buf[682]*(15)+in_buf[683]*(23)+in_buf[684]*(38)+in_buf[685]*(36)+in_buf[686]*(33)+in_buf[687]*(21)+in_buf[688]*(31)+in_buf[689]*(17)+in_buf[690]*(39)+in_buf[691]*(38)+in_buf[692]*(27)+in_buf[693]*(9)+in_buf[694]*(14)+in_buf[695]*(20)+in_buf[696]*(57)+in_buf[697]*(17)+in_buf[698]*(4)+in_buf[699]*(2)+in_buf[700]*(0)+in_buf[701]*(-2)+in_buf[702]*(-22)+in_buf[703]*(-26)+in_buf[704]*(-7)+in_buf[705]*(-7)+in_buf[706]*(11)+in_buf[707]*(6)+in_buf[708]*(9)+in_buf[709]*(8)+in_buf[710]*(5)+in_buf[711]*(-15)+in_buf[712]*(8)+in_buf[713]*(22)+in_buf[714]*(9)+in_buf[715]*(0)+in_buf[716]*(3)+in_buf[717]*(11)+in_buf[718]*(1)+in_buf[719]*(17)+in_buf[720]*(0)+in_buf[721]*(-22)+in_buf[722]*(-13)+in_buf[723]*(11)+in_buf[724]*(39)+in_buf[725]*(-6)+in_buf[726]*(4)+in_buf[727]*(-1)+in_buf[728]*(0)+in_buf[729]*(1)+in_buf[730]*(2)+in_buf[731]*(-5)+in_buf[732]*(10)+in_buf[733]*(24)+in_buf[734]*(3)+in_buf[735]*(-15)+in_buf[736]*(-35)+in_buf[737]*(-46)+in_buf[738]*(-34)+in_buf[739]*(-13)+in_buf[740]*(-9)+in_buf[741]*(-22)+in_buf[742]*(-46)+in_buf[743]*(-41)+in_buf[744]*(-16)+in_buf[745]*(0)+in_buf[746]*(0)+in_buf[747]*(-24)+in_buf[748]*(-46)+in_buf[749]*(-59)+in_buf[750]*(-33)+in_buf[751]*(-3)+in_buf[752]*(0)+in_buf[753]*(-13)+in_buf[754]*(-1)+in_buf[755]*(3)+in_buf[756]*(-3)+in_buf[757]*(-3)+in_buf[758]*(1)+in_buf[759]*(1)+in_buf[760]*(-2)+in_buf[761]*(-20)+in_buf[762]*(-29)+in_buf[763]*(-29)+in_buf[764]*(-44)+in_buf[765]*(-45)+in_buf[766]*(-44)+in_buf[767]*(-19)+in_buf[768]*(-7)+in_buf[769]*(-62)+in_buf[770]*(-63)+in_buf[771]*(-74)+in_buf[772]*(-50)+in_buf[773]*(-40)+in_buf[774]*(-32)+in_buf[775]*(-39)+in_buf[776]*(-42)+in_buf[777]*(-33)+in_buf[778]*(-20)+in_buf[779]*(-16)+in_buf[780]*(-2)+in_buf[781]*(3)+in_buf[782]*(-3)+in_buf[783]*(0);
assign in_buf_weight063=in_buf[0]*(-1)+in_buf[1]*(1)+in_buf[2]*(-2)+in_buf[3]*(0)+in_buf[4]*(0)+in_buf[5]*(4)+in_buf[6]*(-2)+in_buf[7]*(-2)+in_buf[8]*(0)+in_buf[9]*(4)+in_buf[10]*(-2)+in_buf[11]*(2)+in_buf[12]*(11)+in_buf[13]*(4)+in_buf[14]*(-16)+in_buf[15]*(-16)+in_buf[16]*(0)+in_buf[17]*(4)+in_buf[18]*(0)+in_buf[19]*(0)+in_buf[20]*(4)+in_buf[21]*(-3)+in_buf[22]*(2)+in_buf[23]*(-1)+in_buf[24]*(0)+in_buf[25]*(2)+in_buf[26]*(0)+in_buf[27]*(-1)+in_buf[28]*(1)+in_buf[29]*(-3)+in_buf[30]*(0)+in_buf[31]*(4)+in_buf[32]*(6)+in_buf[33]*(5)+in_buf[34]*(-2)+in_buf[35]*(4)+in_buf[36]*(21)+in_buf[37]*(9)+in_buf[38]*(10)+in_buf[39]*(-4)+in_buf[40]*(3)+in_buf[41]*(29)+in_buf[42]*(8)+in_buf[43]*(-16)+in_buf[44]*(-17)+in_buf[45]*(3)+in_buf[46]*(24)+in_buf[47]*(30)+in_buf[48]*(43)+in_buf[49]*(31)+in_buf[50]*(13)+in_buf[51]*(22)+in_buf[52]*(4)+in_buf[53]*(4)+in_buf[54]*(4)+in_buf[55]*(1)+in_buf[56]*(0)+in_buf[57]*(2)+in_buf[58]*(15)+in_buf[59]*(-29)+in_buf[60]*(-18)+in_buf[61]*(9)+in_buf[62]*(17)+in_buf[63]*(36)+in_buf[64]*(19)+in_buf[65]*(-12)+in_buf[66]*(-16)+in_buf[67]*(10)+in_buf[68]*(-5)+in_buf[69]*(-15)+in_buf[70]*(0)+in_buf[71]*(-6)+in_buf[72]*(-12)+in_buf[73]*(6)+in_buf[74]*(19)+in_buf[75]*(11)+in_buf[76]*(10)+in_buf[77]*(11)+in_buf[78]*(30)+in_buf[79]*(-7)+in_buf[80]*(-3)+in_buf[81]*(-13)+in_buf[82]*(2)+in_buf[83]*(3)+in_buf[84]*(-3)+in_buf[85]*(2)+in_buf[86]*(-15)+in_buf[87]*(-32)+in_buf[88]*(-8)+in_buf[89]*(20)+in_buf[90]*(18)+in_buf[91]*(37)+in_buf[92]*(20)+in_buf[93]*(-14)+in_buf[94]*(0)+in_buf[95]*(14)+in_buf[96]*(-11)+in_buf[97]*(-1)+in_buf[98]*(14)+in_buf[99]*(0)+in_buf[100]*(-17)+in_buf[101]*(-13)+in_buf[102]*(-1)+in_buf[103]*(-2)+in_buf[104]*(4)+in_buf[105]*(26)+in_buf[106]*(20)+in_buf[107]*(30)+in_buf[108]*(-1)+in_buf[109]*(-16)+in_buf[110]*(6)+in_buf[111]*(-3)+in_buf[112]*(1)+in_buf[113]*(0)+in_buf[114]*(-18)+in_buf[115]*(-2)+in_buf[116]*(29)+in_buf[117]*(4)+in_buf[118]*(-8)+in_buf[119]*(18)+in_buf[120]*(3)+in_buf[121]*(16)+in_buf[122]*(16)+in_buf[123]*(6)+in_buf[124]*(2)+in_buf[125]*(1)+in_buf[126]*(-4)+in_buf[127]*(-22)+in_buf[128]*(-15)+in_buf[129]*(-7)+in_buf[130]*(-24)+in_buf[131]*(-14)+in_buf[132]*(-1)+in_buf[133]*(7)+in_buf[134]*(10)+in_buf[135]*(35)+in_buf[136]*(28)+in_buf[137]*(2)+in_buf[138]*(-18)+in_buf[139]*(15)+in_buf[140]*(2)+in_buf[141]*(-1)+in_buf[142]*(-15)+in_buf[143]*(-20)+in_buf[144]*(-2)+in_buf[145]*(-20)+in_buf[146]*(-8)+in_buf[147]*(13)+in_buf[148]*(7)+in_buf[149]*(21)+in_buf[150]*(28)+in_buf[151]*(19)+in_buf[152]*(18)+in_buf[153]*(7)+in_buf[154]*(7)+in_buf[155]*(3)+in_buf[156]*(2)+in_buf[157]*(9)+in_buf[158]*(0)+in_buf[159]*(6)+in_buf[160]*(3)+in_buf[161]*(0)+in_buf[162]*(-11)+in_buf[163]*(8)+in_buf[164]*(27)+in_buf[165]*(11)+in_buf[166]*(5)+in_buf[167]*(18)+in_buf[168]*(1)+in_buf[169]*(-17)+in_buf[170]*(-7)+in_buf[171]*(-35)+in_buf[172]*(-29)+in_buf[173]*(-14)+in_buf[174]*(-30)+in_buf[175]*(-6)+in_buf[176]*(7)+in_buf[177]*(8)+in_buf[178]*(4)+in_buf[179]*(-1)+in_buf[180]*(1)+in_buf[181]*(14)+in_buf[182]*(21)+in_buf[183]*(27)+in_buf[184]*(23)+in_buf[185]*(24)+in_buf[186]*(-2)+in_buf[187]*(7)+in_buf[188]*(1)+in_buf[189]*(5)+in_buf[190]*(9)+in_buf[191]*(11)+in_buf[192]*(13)+in_buf[193]*(6)+in_buf[194]*(-5)+in_buf[195]*(-3)+in_buf[196]*(3)+in_buf[197]*(-36)+in_buf[198]*(-1)+in_buf[199]*(-46)+in_buf[200]*(-36)+in_buf[201]*(-7)+in_buf[202]*(-33)+in_buf[203]*(-33)+in_buf[204]*(4)+in_buf[205]*(-1)+in_buf[206]*(-3)+in_buf[207]*(0)+in_buf[208]*(-3)+in_buf[209]*(8)+in_buf[210]*(14)+in_buf[211]*(36)+in_buf[212]*(15)+in_buf[213]*(10)+in_buf[214]*(-2)+in_buf[215]*(-4)+in_buf[216]*(-16)+in_buf[217]*(-2)+in_buf[218]*(0)+in_buf[219]*(14)+in_buf[220]*(17)+in_buf[221]*(-1)+in_buf[222]*(-8)+in_buf[223]*(-18)+in_buf[224]*(-3)+in_buf[225]*(-26)+in_buf[226]*(8)+in_buf[227]*(-2)+in_buf[228]*(-4)+in_buf[229]*(-5)+in_buf[230]*(0)+in_buf[231]*(-22)+in_buf[232]*(6)+in_buf[233]*(-2)+in_buf[234]*(-11)+in_buf[235]*(-6)+in_buf[236]*(-10)+in_buf[237]*(6)+in_buf[238]*(5)+in_buf[239]*(0)+in_buf[240]*(0)+in_buf[241]*(-16)+in_buf[242]*(-11)+in_buf[243]*(-11)+in_buf[244]*(-10)+in_buf[245]*(14)+in_buf[246]*(-12)+in_buf[247]*(-19)+in_buf[248]*(17)+in_buf[249]*(19)+in_buf[250]*(15)+in_buf[251]*(-16)+in_buf[252]*(-7)+in_buf[253]*(-27)+in_buf[254]*(13)+in_buf[255]*(0)+in_buf[256]*(-12)+in_buf[257]*(-19)+in_buf[258]*(-2)+in_buf[259]*(-12)+in_buf[260]*(0)+in_buf[261]*(7)+in_buf[262]*(-4)+in_buf[263]*(0)+in_buf[264]*(-10)+in_buf[265]*(1)+in_buf[266]*(-14)+in_buf[267]*(-26)+in_buf[268]*(-27)+in_buf[269]*(-20)+in_buf[270]*(-23)+in_buf[271]*(-11)+in_buf[272]*(7)+in_buf[273]*(0)+in_buf[274]*(-18)+in_buf[275]*(-8)+in_buf[276]*(12)+in_buf[277]*(-19)+in_buf[278]*(-23)+in_buf[279]*(-27)+in_buf[280]*(-9)+in_buf[281]*(-12)+in_buf[282]*(-17)+in_buf[283]*(0)+in_buf[284]*(-8)+in_buf[285]*(-14)+in_buf[286]*(-19)+in_buf[287]*(-2)+in_buf[288]*(-1)+in_buf[289]*(10)+in_buf[290]*(0)+in_buf[291]*(2)+in_buf[292]*(7)+in_buf[293]*(-10)+in_buf[294]*(-9)+in_buf[295]*(-24)+in_buf[296]*(-30)+in_buf[297]*(-23)+in_buf[298]*(-13)+in_buf[299]*(-9)+in_buf[300]*(-10)+in_buf[301]*(-5)+in_buf[302]*(0)+in_buf[303]*(17)+in_buf[304]*(0)+in_buf[305]*(-33)+in_buf[306]*(-52)+in_buf[307]*(-26)+in_buf[308]*(3)+in_buf[309]*(-28)+in_buf[310]*(-21)+in_buf[311]*(-7)+in_buf[312]*(-22)+in_buf[313]*(-2)+in_buf[314]*(6)+in_buf[315]*(6)+in_buf[316]*(21)+in_buf[317]*(14)+in_buf[318]*(11)+in_buf[319]*(0)+in_buf[320]*(24)+in_buf[321]*(11)+in_buf[322]*(0)+in_buf[323]*(-12)+in_buf[324]*(-1)+in_buf[325]*(7)+in_buf[326]*(-3)+in_buf[327]*(0)+in_buf[328]*(-1)+in_buf[329]*(18)+in_buf[330]*(19)+in_buf[331]*(7)+in_buf[332]*(-2)+in_buf[333]*(-25)+in_buf[334]*(-17)+in_buf[335]*(-45)+in_buf[336]*(-5)+in_buf[337]*(-4)+in_buf[338]*(3)+in_buf[339]*(-9)+in_buf[340]*(-3)+in_buf[341]*(14)+in_buf[342]*(22)+in_buf[343]*(20)+in_buf[344]*(-1)+in_buf[345]*(5)+in_buf[346]*(4)+in_buf[347]*(5)+in_buf[348]*(1)+in_buf[349]*(13)+in_buf[350]*(2)+in_buf[351]*(10)+in_buf[352]*(16)+in_buf[353]*(22)+in_buf[354]*(8)+in_buf[355]*(17)+in_buf[356]*(22)+in_buf[357]*(32)+in_buf[358]*(29)+in_buf[359]*(36)+in_buf[360]*(23)+in_buf[361]*(-32)+in_buf[362]*(-40)+in_buf[363]*(-44)+in_buf[364]*(-15)+in_buf[365]*(2)+in_buf[366]*(-11)+in_buf[367]*(-19)+in_buf[368]*(16)+in_buf[369]*(29)+in_buf[370]*(33)+in_buf[371]*(29)+in_buf[372]*(23)+in_buf[373]*(8)+in_buf[374]*(12)+in_buf[375]*(-3)+in_buf[376]*(-5)+in_buf[377]*(9)+in_buf[378]*(5)+in_buf[379]*(27)+in_buf[380]*(24)+in_buf[381]*(8)+in_buf[382]*(20)+in_buf[383]*(29)+in_buf[384]*(22)+in_buf[385]*(21)+in_buf[386]*(25)+in_buf[387]*(39)+in_buf[388]*(-4)+in_buf[389]*(-17)+in_buf[390]*(-34)+in_buf[391]*(-12)+in_buf[392]*(-11)+in_buf[393]*(-7)+in_buf[394]*(-15)+in_buf[395]*(-10)+in_buf[396]*(6)+in_buf[397]*(34)+in_buf[398]*(26)+in_buf[399]*(33)+in_buf[400]*(24)+in_buf[401]*(14)+in_buf[402]*(9)+in_buf[403]*(6)+in_buf[404]*(10)+in_buf[405]*(8)+in_buf[406]*(3)+in_buf[407]*(14)+in_buf[408]*(18)+in_buf[409]*(10)+in_buf[410]*(17)+in_buf[411]*(28)+in_buf[412]*(28)+in_buf[413]*(29)+in_buf[414]*(15)+in_buf[415]*(7)+in_buf[416]*(-9)+in_buf[417]*(3)+in_buf[418]*(-31)+in_buf[419]*(-16)+in_buf[420]*(-17)+in_buf[421]*(9)+in_buf[422]*(1)+in_buf[423]*(-3)+in_buf[424]*(-10)+in_buf[425]*(-4)+in_buf[426]*(12)+in_buf[427]*(39)+in_buf[428]*(30)+in_buf[429]*(15)+in_buf[430]*(19)+in_buf[431]*(11)+in_buf[432]*(15)+in_buf[433]*(9)+in_buf[434]*(0)+in_buf[435]*(5)+in_buf[436]*(12)+in_buf[437]*(15)+in_buf[438]*(11)+in_buf[439]*(18)+in_buf[440]*(16)+in_buf[441]*(8)+in_buf[442]*(15)+in_buf[443]*(-2)+in_buf[444]*(-22)+in_buf[445]*(14)+in_buf[446]*(-3)+in_buf[447]*(-28)+in_buf[448]*(-2)+in_buf[449]*(4)+in_buf[450]*(-8)+in_buf[451]*(-6)+in_buf[452]*(-16)+in_buf[453]*(-3)+in_buf[454]*(20)+in_buf[455]*(32)+in_buf[456]*(37)+in_buf[457]*(3)+in_buf[458]*(13)+in_buf[459]*(17)+in_buf[460]*(13)+in_buf[461]*(-5)+in_buf[462]*(4)+in_buf[463]*(3)+in_buf[464]*(-1)+in_buf[465]*(11)+in_buf[466]*(22)+in_buf[467]*(-1)+in_buf[468]*(17)+in_buf[469]*(-11)+in_buf[470]*(1)+in_buf[471]*(10)+in_buf[472]*(-4)+in_buf[473]*(9)+in_buf[474]*(-26)+in_buf[475]*(-30)+in_buf[476]*(1)+in_buf[477]*(0)+in_buf[478]*(5)+in_buf[479]*(-12)+in_buf[480]*(-11)+in_buf[481]*(-16)+in_buf[482]*(1)+in_buf[483]*(24)+in_buf[484]*(20)+in_buf[485]*(12)+in_buf[486]*(12)+in_buf[487]*(10)+in_buf[488]*(3)+in_buf[489]*(-4)+in_buf[490]*(-14)+in_buf[491]*(0)+in_buf[492]*(11)+in_buf[493]*(14)+in_buf[494]*(19)+in_buf[495]*(-1)+in_buf[496]*(1)+in_buf[497]*(-4)+in_buf[498]*(-1)+in_buf[499]*(21)+in_buf[500]*(2)+in_buf[501]*(-9)+in_buf[502]*(-14)+in_buf[503]*(-16)+in_buf[504]*(-22)+in_buf[505]*(-7)+in_buf[506]*(-10)+in_buf[507]*(-19)+in_buf[508]*(-14)+in_buf[509]*(-25)+in_buf[510]*(-3)+in_buf[511]*(16)+in_buf[512]*(4)+in_buf[513]*(4)+in_buf[514]*(1)+in_buf[515]*(6)+in_buf[516]*(12)+in_buf[517]*(0)+in_buf[518]*(1)+in_buf[519]*(2)+in_buf[520]*(11)+in_buf[521]*(4)+in_buf[522]*(0)+in_buf[523]*(3)+in_buf[524]*(-4)+in_buf[525]*(-3)+in_buf[526]*(-12)+in_buf[527]*(-10)+in_buf[528]*(-15)+in_buf[529]*(-20)+in_buf[530]*(-39)+in_buf[531]*(-27)+in_buf[532]*(-17)+in_buf[533]*(-20)+in_buf[534]*(-7)+in_buf[535]*(0)+in_buf[536]*(-9)+in_buf[537]*(-8)+in_buf[538]*(-10)+in_buf[539]*(-1)+in_buf[540]*(3)+in_buf[541]*(-5)+in_buf[542]*(3)+in_buf[543]*(0)+in_buf[544]*(-8)+in_buf[545]*(-17)+in_buf[546]*(2)+in_buf[547]*(11)+in_buf[548]*(9)+in_buf[549]*(6)+in_buf[550]*(11)+in_buf[551]*(0)+in_buf[552]*(-11)+in_buf[553]*(-2)+in_buf[554]*(-14)+in_buf[555]*(-15)+in_buf[556]*(-2)+in_buf[557]*(-40)+in_buf[558]*(-11)+in_buf[559]*(-5)+in_buf[560]*(0)+in_buf[561]*(26)+in_buf[562]*(-14)+in_buf[563]*(-29)+in_buf[564]*(-6)+in_buf[565]*(-11)+in_buf[566]*(-16)+in_buf[567]*(-7)+in_buf[568]*(-7)+in_buf[569]*(0)+in_buf[570]*(7)+in_buf[571]*(-13)+in_buf[572]*(-20)+in_buf[573]*(-6)+in_buf[574]*(9)+in_buf[575]*(8)+in_buf[576]*(2)+in_buf[577]*(0)+in_buf[578]*(9)+in_buf[579]*(-9)+in_buf[580]*(-5)+in_buf[581]*(-7)+in_buf[582]*(-10)+in_buf[583]*(-26)+in_buf[584]*(5)+in_buf[585]*(-17)+in_buf[586]*(-18)+in_buf[587]*(2)+in_buf[588]*(-20)+in_buf[589]*(-18)+in_buf[590]*(-33)+in_buf[591]*(-39)+in_buf[592]*(-5)+in_buf[593]*(-15)+in_buf[594]*(-7)+in_buf[595]*(-2)+in_buf[596]*(7)+in_buf[597]*(4)+in_buf[598]*(-9)+in_buf[599]*(3)+in_buf[600]*(-1)+in_buf[601]*(10)+in_buf[602]*(12)+in_buf[603]*(5)+in_buf[604]*(10)+in_buf[605]*(17)+in_buf[606]*(-8)+in_buf[607]*(-3)+in_buf[608]*(-16)+in_buf[609]*(-21)+in_buf[610]*(-11)+in_buf[611]*(-13)+in_buf[612]*(-21)+in_buf[613]*(-36)+in_buf[614]*(-21)+in_buf[615]*(6)+in_buf[616]*(-21)+in_buf[617]*(-12)+in_buf[618]*(-31)+in_buf[619]*(-13)+in_buf[620]*(-10)+in_buf[621]*(-30)+in_buf[622]*(0)+in_buf[623]*(0)+in_buf[624]*(-6)+in_buf[625]*(-7)+in_buf[626]*(3)+in_buf[627]*(16)+in_buf[628]*(16)+in_buf[629]*(14)+in_buf[630]*(11)+in_buf[631]*(6)+in_buf[632]*(9)+in_buf[633]*(1)+in_buf[634]*(-4)+in_buf[635]*(-7)+in_buf[636]*(-24)+in_buf[637]*(-15)+in_buf[638]*(13)+in_buf[639]*(10)+in_buf[640]*(-17)+in_buf[641]*(-24)+in_buf[642]*(-2)+in_buf[643]*(1)+in_buf[644]*(0)+in_buf[645]*(1)+in_buf[646]*(-23)+in_buf[647]*(5)+in_buf[648]*(-1)+in_buf[649]*(-16)+in_buf[650]*(-15)+in_buf[651]*(-2)+in_buf[652]*(17)+in_buf[653]*(-1)+in_buf[654]*(9)+in_buf[655]*(-2)+in_buf[656]*(-2)+in_buf[657]*(0)+in_buf[658]*(4)+in_buf[659]*(4)+in_buf[660]*(6)+in_buf[661]*(0)+in_buf[662]*(10)+in_buf[663]*(1)+in_buf[664]*(-6)+in_buf[665]*(21)+in_buf[666]*(8)+in_buf[667]*(-6)+in_buf[668]*(-15)+in_buf[669]*(-27)+in_buf[670]*(-27)+in_buf[671]*(-2)+in_buf[672]*(3)+in_buf[673]*(4)+in_buf[674]*(-23)+in_buf[675]*(-10)+in_buf[676]*(-11)+in_buf[677]*(-3)+in_buf[678]*(-1)+in_buf[679]*(13)+in_buf[680]*(12)+in_buf[681]*(14)+in_buf[682]*(17)+in_buf[683]*(12)+in_buf[684]*(14)+in_buf[685]*(12)+in_buf[686]*(-1)+in_buf[687]*(3)+in_buf[688]*(11)+in_buf[689]*(-16)+in_buf[690]*(-11)+in_buf[691]*(0)+in_buf[692]*(16)+in_buf[693]*(-7)+in_buf[694]*(21)+in_buf[695]*(19)+in_buf[696]*(-38)+in_buf[697]*(-9)+in_buf[698]*(-18)+in_buf[699]*(1)+in_buf[700]*(-2)+in_buf[701]*(1)+in_buf[702]*(32)+in_buf[703]*(-6)+in_buf[704]*(-14)+in_buf[705]*(-4)+in_buf[706]*(-17)+in_buf[707]*(-8)+in_buf[708]*(-10)+in_buf[709]*(-2)+in_buf[710]*(11)+in_buf[711]*(5)+in_buf[712]*(-21)+in_buf[713]*(-13)+in_buf[714]*(-10)+in_buf[715]*(-10)+in_buf[716]*(-19)+in_buf[717]*(-22)+in_buf[718]*(3)+in_buf[719]*(2)+in_buf[720]*(1)+in_buf[721]*(0)+in_buf[722]*(-5)+in_buf[723]*(-17)+in_buf[724]*(-29)+in_buf[725]*(7)+in_buf[726]*(-8)+in_buf[727]*(-2)+in_buf[728]*(0)+in_buf[729]*(0)+in_buf[730]*(3)+in_buf[731]*(6)+in_buf[732]*(39)+in_buf[733]*(39)+in_buf[734]*(35)+in_buf[735]*(17)+in_buf[736]*(0)+in_buf[737]*(-13)+in_buf[738]*(-4)+in_buf[739]*(2)+in_buf[740]*(15)+in_buf[741]*(-2)+in_buf[742]*(15)+in_buf[743]*(-1)+in_buf[744]*(8)+in_buf[745]*(1)+in_buf[746]*(-2)+in_buf[747]*(-19)+in_buf[748]*(-10)+in_buf[749]*(-13)+in_buf[750]*(-6)+in_buf[751]*(13)+in_buf[752]*(24)+in_buf[753]*(1)+in_buf[754]*(3)+in_buf[755]*(-1)+in_buf[756]*(1)+in_buf[757]*(1)+in_buf[758]*(-2)+in_buf[759]*(-3)+in_buf[760]*(-21)+in_buf[761]*(-22)+in_buf[762]*(-12)+in_buf[763]*(-4)+in_buf[764]*(-7)+in_buf[765]*(-15)+in_buf[766]*(-16)+in_buf[767]*(3)+in_buf[768]*(2)+in_buf[769]*(-37)+in_buf[770]*(-14)+in_buf[771]*(14)+in_buf[772]*(-10)+in_buf[773]*(-23)+in_buf[774]*(-5)+in_buf[775]*(21)+in_buf[776]*(7)+in_buf[777]*(-17)+in_buf[778]*(-31)+in_buf[779]*(-25)+in_buf[780]*(2)+in_buf[781]*(-2)+in_buf[782]*(4)+in_buf[783]*(4);
wire [DATAWIDTH-1:0]   weight0_bias00;
wire [DATAWIDTH-1:0]   weight0_bias01;
wire [DATAWIDTH-1:0]   weight0_bias02;
wire [DATAWIDTH-1:0]   weight0_bias03;
wire [DATAWIDTH-1:0]   weight0_bias04;
wire [DATAWIDTH-1:0]   weight0_bias05;
wire [DATAWIDTH-1:0]   weight0_bias06;
wire [DATAWIDTH-1:0]   weight0_bias07;
wire [DATAWIDTH-1:0]   weight0_bias08;
wire [DATAWIDTH-1:0]   weight0_bias09;
wire [DATAWIDTH-1:0]   weight0_bias010;
wire [DATAWIDTH-1:0]   weight0_bias011;
wire [DATAWIDTH-1:0]   weight0_bias012;
wire [DATAWIDTH-1:0]   weight0_bias013;
wire [DATAWIDTH-1:0]   weight0_bias014;
wire [DATAWIDTH-1:0]   weight0_bias015;
wire [DATAWIDTH-1:0]   weight0_bias016;
wire [DATAWIDTH-1:0]   weight0_bias017;
wire [DATAWIDTH-1:0]   weight0_bias018;
wire [DATAWIDTH-1:0]   weight0_bias019;
wire [DATAWIDTH-1:0]   weight0_bias020;
wire [DATAWIDTH-1:0]   weight0_bias021;
wire [DATAWIDTH-1:0]   weight0_bias022;
wire [DATAWIDTH-1:0]   weight0_bias023;
wire [DATAWIDTH-1:0]   weight0_bias024;
wire [DATAWIDTH-1:0]   weight0_bias025;
wire [DATAWIDTH-1:0]   weight0_bias026;
wire [DATAWIDTH-1:0]   weight0_bias027;
wire [DATAWIDTH-1:0]   weight0_bias028;
wire [DATAWIDTH-1:0]   weight0_bias029;
wire [DATAWIDTH-1:0]   weight0_bias030;
wire [DATAWIDTH-1:0]   weight0_bias031;
wire [DATAWIDTH-1:0]   weight0_bias032;
wire [DATAWIDTH-1:0]   weight0_bias033;
wire [DATAWIDTH-1:0]   weight0_bias034;
wire [DATAWIDTH-1:0]   weight0_bias035;
wire [DATAWIDTH-1:0]   weight0_bias036;
wire [DATAWIDTH-1:0]   weight0_bias037;
wire [DATAWIDTH-1:0]   weight0_bias038;
wire [DATAWIDTH-1:0]   weight0_bias039;
wire [DATAWIDTH-1:0]   weight0_bias040;
wire [DATAWIDTH-1:0]   weight0_bias041;
wire [DATAWIDTH-1:0]   weight0_bias042;
wire [DATAWIDTH-1:0]   weight0_bias043;
wire [DATAWIDTH-1:0]   weight0_bias044;
wire [DATAWIDTH-1:0]   weight0_bias045;
wire [DATAWIDTH-1:0]   weight0_bias046;
wire [DATAWIDTH-1:0]   weight0_bias047;
wire [DATAWIDTH-1:0]   weight0_bias048;
wire [DATAWIDTH-1:0]   weight0_bias049;
wire [DATAWIDTH-1:0]   weight0_bias050;
wire [DATAWIDTH-1:0]   weight0_bias051;
wire [DATAWIDTH-1:0]   weight0_bias052;
wire [DATAWIDTH-1:0]   weight0_bias053;
wire [DATAWIDTH-1:0]   weight0_bias054;
wire [DATAWIDTH-1:0]   weight0_bias055;
wire [DATAWIDTH-1:0]   weight0_bias056;
wire [DATAWIDTH-1:0]   weight0_bias057;
wire [DATAWIDTH-1:0]   weight0_bias058;
wire [DATAWIDTH-1:0]   weight0_bias059;
wire [DATAWIDTH-1:0]   weight0_bias060;
wire [DATAWIDTH-1:0]   weight0_bias061;
wire [DATAWIDTH-1:0]   weight0_bias062;
wire [DATAWIDTH-1:0]   weight0_bias063;
assign weight0_bias00=in_buf_weight00+(22);
assign weight0_bias01=in_buf_weight01+(0);
assign weight0_bias02=in_buf_weight02+(7);
assign weight0_bias03=in_buf_weight03+(-4);
assign weight0_bias04=in_buf_weight04+(11);
assign weight0_bias05=in_buf_weight05+(6);
assign weight0_bias06=in_buf_weight06+(3);
assign weight0_bias07=in_buf_weight07+(24);
assign weight0_bias08=in_buf_weight08+(3);
assign weight0_bias09=in_buf_weight09+(-5);
assign weight0_bias010=in_buf_weight010+(-8);
assign weight0_bias011=in_buf_weight011+(-1);
assign weight0_bias012=in_buf_weight012+(-1);
assign weight0_bias013=in_buf_weight013+(22);
assign weight0_bias014=in_buf_weight014+(0);
assign weight0_bias015=in_buf_weight015+(28);
assign weight0_bias016=in_buf_weight016+(17);
assign weight0_bias017=in_buf_weight017+(3);
assign weight0_bias018=in_buf_weight018+(14);
assign weight0_bias019=in_buf_weight019+(28);
assign weight0_bias020=in_buf_weight020+(12);
assign weight0_bias021=in_buf_weight021+(17);
assign weight0_bias022=in_buf_weight022+(21);
assign weight0_bias023=in_buf_weight023+(16);
assign weight0_bias024=in_buf_weight024+(1);
assign weight0_bias025=in_buf_weight025+(10);
assign weight0_bias026=in_buf_weight026+(3);
assign weight0_bias027=in_buf_weight027+(-3);
assign weight0_bias028=in_buf_weight028+(43);
assign weight0_bias029=in_buf_weight029+(32);
assign weight0_bias030=in_buf_weight030+(-4);
assign weight0_bias031=in_buf_weight031+(-2);
assign weight0_bias032=in_buf_weight032+(19);
assign weight0_bias033=in_buf_weight033+(51);
assign weight0_bias034=in_buf_weight034+(22);
assign weight0_bias035=in_buf_weight035+(29);
assign weight0_bias036=in_buf_weight036+(3);
assign weight0_bias037=in_buf_weight037+(12);
assign weight0_bias038=in_buf_weight038+(-4);
assign weight0_bias039=in_buf_weight039+(5);
assign weight0_bias040=in_buf_weight040+(-12);
assign weight0_bias041=in_buf_weight041+(18);
assign weight0_bias042=in_buf_weight042+(4);
assign weight0_bias043=in_buf_weight043+(2);
assign weight0_bias044=in_buf_weight044+(-2);
assign weight0_bias045=in_buf_weight045+(13);
assign weight0_bias046=in_buf_weight046+(14);
assign weight0_bias047=in_buf_weight047+(-21);
assign weight0_bias048=in_buf_weight048+(3);
assign weight0_bias049=in_buf_weight049+(8);
assign weight0_bias050=in_buf_weight050+(14);
assign weight0_bias051=in_buf_weight051+(-2);
assign weight0_bias052=in_buf_weight052+(6);
assign weight0_bias053=in_buf_weight053+(-3);
assign weight0_bias054=in_buf_weight054+(-2);
assign weight0_bias055=in_buf_weight055+(18);
assign weight0_bias056=in_buf_weight056+(-4);
assign weight0_bias057=in_buf_weight057+(20);
assign weight0_bias058=in_buf_weight058+(-10);
assign weight0_bias059=in_buf_weight059+(11);
assign weight0_bias060=in_buf_weight060+(38);
assign weight0_bias061=in_buf_weight061+(-1);
assign weight0_bias062=in_buf_weight062+(-7);
assign weight0_bias063=in_buf_weight063+(1);
wire [DATAWIDTH-1:0]   bias0_relu00;
wire [DATAWIDTH-1:0]   bias0_relu01;
wire [DATAWIDTH-1:0]   bias0_relu02;
wire [DATAWIDTH-1:0]   bias0_relu03;
wire [DATAWIDTH-1:0]   bias0_relu04;
wire [DATAWIDTH-1:0]   bias0_relu05;
wire [DATAWIDTH-1:0]   bias0_relu06;
wire [DATAWIDTH-1:0]   bias0_relu07;
wire [DATAWIDTH-1:0]   bias0_relu08;
wire [DATAWIDTH-1:0]   bias0_relu09;
wire [DATAWIDTH-1:0]   bias0_relu010;
wire [DATAWIDTH-1:0]   bias0_relu011;
wire [DATAWIDTH-1:0]   bias0_relu012;
wire [DATAWIDTH-1:0]   bias0_relu013;
wire [DATAWIDTH-1:0]   bias0_relu014;
wire [DATAWIDTH-1:0]   bias0_relu015;
wire [DATAWIDTH-1:0]   bias0_relu016;
wire [DATAWIDTH-1:0]   bias0_relu017;
wire [DATAWIDTH-1:0]   bias0_relu018;
wire [DATAWIDTH-1:0]   bias0_relu019;
wire [DATAWIDTH-1:0]   bias0_relu020;
wire [DATAWIDTH-1:0]   bias0_relu021;
wire [DATAWIDTH-1:0]   bias0_relu022;
wire [DATAWIDTH-1:0]   bias0_relu023;
wire [DATAWIDTH-1:0]   bias0_relu024;
wire [DATAWIDTH-1:0]   bias0_relu025;
wire [DATAWIDTH-1:0]   bias0_relu026;
wire [DATAWIDTH-1:0]   bias0_relu027;
wire [DATAWIDTH-1:0]   bias0_relu028;
wire [DATAWIDTH-1:0]   bias0_relu029;
wire [DATAWIDTH-1:0]   bias0_relu030;
wire [DATAWIDTH-1:0]   bias0_relu031;
wire [DATAWIDTH-1:0]   bias0_relu032;
wire [DATAWIDTH-1:0]   bias0_relu033;
wire [DATAWIDTH-1:0]   bias0_relu034;
wire [DATAWIDTH-1:0]   bias0_relu035;
wire [DATAWIDTH-1:0]   bias0_relu036;
wire [DATAWIDTH-1:0]   bias0_relu037;
wire [DATAWIDTH-1:0]   bias0_relu038;
wire [DATAWIDTH-1:0]   bias0_relu039;
wire [DATAWIDTH-1:0]   bias0_relu040;
wire [DATAWIDTH-1:0]   bias0_relu041;
wire [DATAWIDTH-1:0]   bias0_relu042;
wire [DATAWIDTH-1:0]   bias0_relu043;
wire [DATAWIDTH-1:0]   bias0_relu044;
wire [DATAWIDTH-1:0]   bias0_relu045;
wire [DATAWIDTH-1:0]   bias0_relu046;
wire [DATAWIDTH-1:0]   bias0_relu047;
wire [DATAWIDTH-1:0]   bias0_relu048;
wire [DATAWIDTH-1:0]   bias0_relu049;
wire [DATAWIDTH-1:0]   bias0_relu050;
wire [DATAWIDTH-1:0]   bias0_relu051;
wire [DATAWIDTH-1:0]   bias0_relu052;
wire [DATAWIDTH-1:0]   bias0_relu053;
wire [DATAWIDTH-1:0]   bias0_relu054;
wire [DATAWIDTH-1:0]   bias0_relu055;
wire [DATAWIDTH-1:0]   bias0_relu056;
wire [DATAWIDTH-1:0]   bias0_relu057;
wire [DATAWIDTH-1:0]   bias0_relu058;
wire [DATAWIDTH-1:0]   bias0_relu059;
wire [DATAWIDTH-1:0]   bias0_relu060;
wire [DATAWIDTH-1:0]   bias0_relu061;
wire [DATAWIDTH-1:0]   bias0_relu062;
wire [DATAWIDTH-1:0]   bias0_relu063;
assign bias0_relu00=(weight0_bias00[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias00;
assign bias0_relu01=(weight0_bias01[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias01;
assign bias0_relu02=(weight0_bias02[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias02;
assign bias0_relu03=(weight0_bias03[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias03;
assign bias0_relu04=(weight0_bias04[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias04;
assign bias0_relu05=(weight0_bias05[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias05;
assign bias0_relu06=(weight0_bias06[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias06;
assign bias0_relu07=(weight0_bias07[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias07;
assign bias0_relu08=(weight0_bias08[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias08;
assign bias0_relu09=(weight0_bias09[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias09;
assign bias0_relu010=(weight0_bias010[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias010;
assign bias0_relu011=(weight0_bias011[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias011;
assign bias0_relu012=(weight0_bias012[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias012;
assign bias0_relu013=(weight0_bias013[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias013;
assign bias0_relu014=(weight0_bias014[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias014;
assign bias0_relu015=(weight0_bias015[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias015;
assign bias0_relu016=(weight0_bias016[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias016;
assign bias0_relu017=(weight0_bias017[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias017;
assign bias0_relu018=(weight0_bias018[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias018;
assign bias0_relu019=(weight0_bias019[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias019;
assign bias0_relu020=(weight0_bias020[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias020;
assign bias0_relu021=(weight0_bias021[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias021;
assign bias0_relu022=(weight0_bias022[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias022;
assign bias0_relu023=(weight0_bias023[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias023;
assign bias0_relu024=(weight0_bias024[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias024;
assign bias0_relu025=(weight0_bias025[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias025;
assign bias0_relu026=(weight0_bias026[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias026;
assign bias0_relu027=(weight0_bias027[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias027;
assign bias0_relu028=(weight0_bias028[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias028;
assign bias0_relu029=(weight0_bias029[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias029;
assign bias0_relu030=(weight0_bias030[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias030;
assign bias0_relu031=(weight0_bias031[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias031;
assign bias0_relu032=(weight0_bias032[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias032;
assign bias0_relu033=(weight0_bias033[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias033;
assign bias0_relu034=(weight0_bias034[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias034;
assign bias0_relu035=(weight0_bias035[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias035;
assign bias0_relu036=(weight0_bias036[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias036;
assign bias0_relu037=(weight0_bias037[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias037;
assign bias0_relu038=(weight0_bias038[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias038;
assign bias0_relu039=(weight0_bias039[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias039;
assign bias0_relu040=(weight0_bias040[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias040;
assign bias0_relu041=(weight0_bias041[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias041;
assign bias0_relu042=(weight0_bias042[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias042;
assign bias0_relu043=(weight0_bias043[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias043;
assign bias0_relu044=(weight0_bias044[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias044;
assign bias0_relu045=(weight0_bias045[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias045;
assign bias0_relu046=(weight0_bias046[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias046;
assign bias0_relu047=(weight0_bias047[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias047;
assign bias0_relu048=(weight0_bias048[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias048;
assign bias0_relu049=(weight0_bias049[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias049;
assign bias0_relu050=(weight0_bias050[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias050;
assign bias0_relu051=(weight0_bias051[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias051;
assign bias0_relu052=(weight0_bias052[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias052;
assign bias0_relu053=(weight0_bias053[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias053;
assign bias0_relu054=(weight0_bias054[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias054;
assign bias0_relu055=(weight0_bias055[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias055;
assign bias0_relu056=(weight0_bias056[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias056;
assign bias0_relu057=(weight0_bias057[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias057;
assign bias0_relu058=(weight0_bias058[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias058;
assign bias0_relu059=(weight0_bias059[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias059;
assign bias0_relu060=(weight0_bias060[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias060;
assign bias0_relu061=(weight0_bias061[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias061;
assign bias0_relu062=(weight0_bias062[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias062;
assign bias0_relu063=(weight0_bias063[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight0_bias063;

wire [DATAWIDTH-1:0]   relu0_weight20;
wire [DATAWIDTH-1:0]   relu0_weight21;
wire [DATAWIDTH-1:0]   relu0_weight22;
wire [DATAWIDTH-1:0]   relu0_weight23;
wire [DATAWIDTH-1:0]   relu0_weight24;
wire [DATAWIDTH-1:0]   relu0_weight25;
wire [DATAWIDTH-1:0]   relu0_weight26;
wire [DATAWIDTH-1:0]   relu0_weight27;
wire [DATAWIDTH-1:0]   relu0_weight28;
wire [DATAWIDTH-1:0]   relu0_weight29;
wire [DATAWIDTH-1:0]   relu0_weight210;
wire [DATAWIDTH-1:0]   relu0_weight211;
wire [DATAWIDTH-1:0]   relu0_weight212;
wire [DATAWIDTH-1:0]   relu0_weight213;
wire [DATAWIDTH-1:0]   relu0_weight214;
wire [DATAWIDTH-1:0]   relu0_weight215;
wire [DATAWIDTH-1:0]   relu0_weight216;
wire [DATAWIDTH-1:0]   relu0_weight217;
wire [DATAWIDTH-1:0]   relu0_weight218;
wire [DATAWIDTH-1:0]   relu0_weight219;
wire [DATAWIDTH-1:0]   relu0_weight220;
wire [DATAWIDTH-1:0]   relu0_weight221;
wire [DATAWIDTH-1:0]   relu0_weight222;
wire [DATAWIDTH-1:0]   relu0_weight223;
wire [DATAWIDTH-1:0]   relu0_weight224;
wire [DATAWIDTH-1:0]   relu0_weight225;
wire [DATAWIDTH-1:0]   relu0_weight226;
wire [DATAWIDTH-1:0]   relu0_weight227;
wire [DATAWIDTH-1:0]   relu0_weight228;
wire [DATAWIDTH-1:0]   relu0_weight229;
wire [DATAWIDTH-1:0]   relu0_weight230;
wire [DATAWIDTH-1:0]   relu0_weight231;
assign relu0_weight20=bias0_relu00*(-8)+bias0_relu01*(-11)+bias0_relu02*(8)+bias0_relu03*(35)+bias0_relu04*(-16)+bias0_relu05*(17)+bias0_relu06*(5)+bias0_relu07*(7)+bias0_relu08*(24)+bias0_relu09*(-2)+bias0_relu010*(-5)+bias0_relu011*(7)+bias0_relu012*(-12)+bias0_relu013*(9)+bias0_relu014*(2)+bias0_relu015*(-28)+bias0_relu016*(72)+bias0_relu017*(22)+bias0_relu018*(-28)+bias0_relu019*(-12)+bias0_relu020*(25)+bias0_relu021*(46)+bias0_relu022*(14)+bias0_relu023*(-16)+bias0_relu024*(10)+bias0_relu025*(-15)+bias0_relu026*(18)+bias0_relu027*(-2)+bias0_relu028*(-37)+bias0_relu029*(16)+bias0_relu030*(38)+bias0_relu031*(5)+bias0_relu032*(-31)+bias0_relu033*(4)+bias0_relu034*(-26)+bias0_relu035*(8)+bias0_relu036*(21)+bias0_relu037*(21)+bias0_relu038*(-7)+bias0_relu039*(-18)+bias0_relu040*(34)+bias0_relu041*(-29)+bias0_relu042*(0)+bias0_relu043*(0)+bias0_relu044*(-25)+bias0_relu045*(-38)+bias0_relu046*(-8)+bias0_relu047*(-27)+bias0_relu048*(-2)+bias0_relu049*(-5)+bias0_relu050*(8)+bias0_relu051*(31)+bias0_relu052*(-9)+bias0_relu053*(3)+bias0_relu054*(25)+bias0_relu055*(1)+bias0_relu056*(2)+bias0_relu057*(37)+bias0_relu058*(26)+bias0_relu059*(-7)+bias0_relu060*(-12)+bias0_relu061*(9)+bias0_relu062*(-13)+bias0_relu063*(22);
assign relu0_weight21=bias0_relu00*(20)+bias0_relu01*(-29)+bias0_relu02*(49)+bias0_relu03*(14)+bias0_relu04*(-1)+bias0_relu05*(28)+bias0_relu06*(-11)+bias0_relu07*(0)+bias0_relu08*(24)+bias0_relu09*(12)+bias0_relu010*(-16)+bias0_relu011*(-3)+bias0_relu012*(36)+bias0_relu013*(16)+bias0_relu014*(-3)+bias0_relu015*(-11)+bias0_relu016*(-16)+bias0_relu017*(32)+bias0_relu018*(-7)+bias0_relu019*(36)+bias0_relu020*(-28)+bias0_relu021*(28)+bias0_relu022*(-46)+bias0_relu023*(-2)+bias0_relu024*(-14)+bias0_relu025*(-20)+bias0_relu026*(40)+bias0_relu027*(-1)+bias0_relu028*(-9)+bias0_relu029*(16)+bias0_relu030*(-11)+bias0_relu031*(-54)+bias0_relu032*(7)+bias0_relu033*(21)+bias0_relu034*(6)+bias0_relu035*(-10)+bias0_relu036*(-64)+bias0_relu037*(33)+bias0_relu038*(12)+bias0_relu039*(22)+bias0_relu040*(11)+bias0_relu041*(5)+bias0_relu042*(38)+bias0_relu043*(26)+bias0_relu044*(8)+bias0_relu045*(3)+bias0_relu046*(45)+bias0_relu047*(-55)+bias0_relu048*(-15)+bias0_relu049*(9)+bias0_relu050*(17)+bias0_relu051*(-40)+bias0_relu052*(-5)+bias0_relu053*(23)+bias0_relu054*(25)+bias0_relu055*(1)+bias0_relu056*(-9)+bias0_relu057*(13)+bias0_relu058*(8)+bias0_relu059*(-26)+bias0_relu060*(59)+bias0_relu061*(-52)+bias0_relu062*(28)+bias0_relu063*(-17);
assign relu0_weight22=bias0_relu00*(-52)+bias0_relu01*(-6)+bias0_relu02*(-10)+bias0_relu03*(55)+bias0_relu04*(3)+bias0_relu05*(34)+bias0_relu06*(15)+bias0_relu07*(20)+bias0_relu08*(13)+bias0_relu09*(0)+bias0_relu010*(22)+bias0_relu011*(45)+bias0_relu012*(57)+bias0_relu013*(-22)+bias0_relu014*(26)+bias0_relu015*(-44)+bias0_relu016*(8)+bias0_relu017*(38)+bias0_relu018*(-14)+bias0_relu019*(-4)+bias0_relu020*(-35)+bias0_relu021*(-13)+bias0_relu022*(-16)+bias0_relu023*(-17)+bias0_relu024*(23)+bias0_relu025*(-23)+bias0_relu026*(4)+bias0_relu027*(-9)+bias0_relu028*(-33)+bias0_relu029*(45)+bias0_relu030*(3)+bias0_relu031*(-32)+bias0_relu032*(39)+bias0_relu033*(17)+bias0_relu034*(9)+bias0_relu035*(-26)+bias0_relu036*(-7)+bias0_relu037*(17)+bias0_relu038*(37)+bias0_relu039*(-2)+bias0_relu040*(35)+bias0_relu041*(-27)+bias0_relu042*(19)+bias0_relu043*(44)+bias0_relu044*(-36)+bias0_relu045*(-10)+bias0_relu046*(10)+bias0_relu047*(15)+bias0_relu048*(20)+bias0_relu049*(35)+bias0_relu050*(12)+bias0_relu051*(-14)+bias0_relu052*(7)+bias0_relu053*(2)+bias0_relu054*(22)+bias0_relu055*(23)+bias0_relu056*(9)+bias0_relu057*(-6)+bias0_relu058*(23)+bias0_relu059*(-51)+bias0_relu060*(21)+bias0_relu061*(-30)+bias0_relu062*(48)+bias0_relu063*(13);
assign relu0_weight23=bias0_relu00*(-57)+bias0_relu01*(-37)+bias0_relu02*(4)+bias0_relu03*(-31)+bias0_relu04*(8)+bias0_relu05*(13)+bias0_relu06*(-12)+bias0_relu07*(16)+bias0_relu08*(11)+bias0_relu09*(7)+bias0_relu010*(46)+bias0_relu011*(11)+bias0_relu012*(19)+bias0_relu013*(-75)+bias0_relu014*(-17)+bias0_relu015*(-2)+bias0_relu016*(-10)+bias0_relu017*(43)+bias0_relu018*(-7)+bias0_relu019*(24)+bias0_relu020*(13)+bias0_relu021*(-42)+bias0_relu022*(17)+bias0_relu023*(16)+bias0_relu024*(18)+bias0_relu025*(7)+bias0_relu026*(-10)+bias0_relu027*(-7)+bias0_relu028*(0)+bias0_relu029*(8)+bias0_relu030*(-1)+bias0_relu031*(-13)+bias0_relu032*(22)+bias0_relu033*(0)+bias0_relu034*(18)+bias0_relu035*(1)+bias0_relu036*(-9)+bias0_relu037*(16)+bias0_relu038*(-1)+bias0_relu039*(28)+bias0_relu040*(56)+bias0_relu041*(18)+bias0_relu042*(22)+bias0_relu043*(16)+bias0_relu044*(0)+bias0_relu045*(-48)+bias0_relu046*(20)+bias0_relu047*(-30)+bias0_relu048*(21)+bias0_relu049*(9)+bias0_relu050*(-9)+bias0_relu051*(-2)+bias0_relu052*(-57)+bias0_relu053*(30)+bias0_relu054*(41)+bias0_relu055*(34)+bias0_relu056*(-11)+bias0_relu057*(29)+bias0_relu058*(35)+bias0_relu059*(-22)+bias0_relu060*(-38)+bias0_relu061*(-13)+bias0_relu062*(-28)+bias0_relu063*(21);
assign relu0_weight24=bias0_relu00*(-26)+bias0_relu01*(17)+bias0_relu02*(47)+bias0_relu03*(14)+bias0_relu04*(0)+bias0_relu05*(35)+bias0_relu06*(-12)+bias0_relu07*(-1)+bias0_relu08*(12)+bias0_relu09*(-4)+bias0_relu010*(-7)+bias0_relu011*(28)+bias0_relu012*(3)+bias0_relu013*(41)+bias0_relu014*(24)+bias0_relu015*(-13)+bias0_relu016*(7)+bias0_relu017*(14)+bias0_relu018*(-20)+bias0_relu019*(34)+bias0_relu020*(-3)+bias0_relu021*(22)+bias0_relu022*(-49)+bias0_relu023*(-15)+bias0_relu024*(13)+bias0_relu025*(-45)+bias0_relu026*(7)+bias0_relu027*(-8)+bias0_relu028*(-30)+bias0_relu029*(-1)+bias0_relu030*(35)+bias0_relu031*(-1)+bias0_relu032*(-3)+bias0_relu033*(17)+bias0_relu034*(2)+bias0_relu035*(21)+bias0_relu036*(-74)+bias0_relu037*(-14)+bias0_relu038*(-5)+bias0_relu039*(17)+bias0_relu040*(-3)+bias0_relu041*(-4)+bias0_relu042*(-15)+bias0_relu043*(27)+bias0_relu044*(15)+bias0_relu045*(15)+bias0_relu046*(12)+bias0_relu047*(-75)+bias0_relu048*(10)+bias0_relu049*(42)+bias0_relu050*(45)+bias0_relu051*(15)+bias0_relu052*(-40)+bias0_relu053*(32)+bias0_relu054*(5)+bias0_relu055*(-7)+bias0_relu056*(15)+bias0_relu057*(4)+bias0_relu058*(31)+bias0_relu059*(-12)+bias0_relu060*(50)+bias0_relu061*(-1)+bias0_relu062*(37)+bias0_relu063*(11);
assign relu0_weight25=bias0_relu00*(-24)+bias0_relu01*(-43)+bias0_relu02*(0)+bias0_relu03*(-12)+bias0_relu04*(16)+bias0_relu05*(3)+bias0_relu06*(-5)+bias0_relu07*(20)+bias0_relu08*(-6)+bias0_relu09*(3)+bias0_relu010*(43)+bias0_relu011*(1)+bias0_relu012*(6)+bias0_relu013*(-65)+bias0_relu014*(-10)+bias0_relu015*(39)+bias0_relu016*(-35)+bias0_relu017*(-1)+bias0_relu018*(16)+bias0_relu019*(31)+bias0_relu020*(11)+bias0_relu021*(5)+bias0_relu022*(22)+bias0_relu023*(-8)+bias0_relu024*(31)+bias0_relu025*(10)+bias0_relu026*(-6)+bias0_relu027*(1)+bias0_relu028*(40)+bias0_relu029*(1)+bias0_relu030*(-10)+bias0_relu031*(-43)+bias0_relu032*(51)+bias0_relu033*(17)+bias0_relu034*(25)+bias0_relu035*(-29)+bias0_relu036*(50)+bias0_relu037*(57)+bias0_relu038*(3)+bias0_relu039*(30)+bias0_relu040*(22)+bias0_relu041*(30)+bias0_relu042*(31)+bias0_relu043*(19)+bias0_relu044*(-17)+bias0_relu045*(-9)+bias0_relu046*(-6)+bias0_relu047*(52)+bias0_relu048*(-4)+bias0_relu049*(1)+bias0_relu050*(12)+bias0_relu051*(-20)+bias0_relu052*(-33)+bias0_relu053*(-24)+bias0_relu054*(-4)+bias0_relu055*(42)+bias0_relu056*(2)+bias0_relu057*(-3)+bias0_relu058*(-9)+bias0_relu059*(8)+bias0_relu060*(15)+bias0_relu061*(-36)+bias0_relu062*(-22)+bias0_relu063*(1);
assign relu0_weight26=bias0_relu00*(12)+bias0_relu01*(-7)+bias0_relu02*(-68)+bias0_relu03*(-14)+bias0_relu04*(34)+bias0_relu05*(24)+bias0_relu06*(6)+bias0_relu07*(22)+bias0_relu08*(0)+bias0_relu09*(5)+bias0_relu010*(42)+bias0_relu011*(22)+bias0_relu012*(-10)+bias0_relu013*(-74)+bias0_relu014*(12)+bias0_relu015*(11)+bias0_relu016*(24)+bias0_relu017*(-7)+bias0_relu018*(60)+bias0_relu019*(-42)+bias0_relu020*(-14)+bias0_relu021*(-40)+bias0_relu022*(21)+bias0_relu023*(47)+bias0_relu024*(4)+bias0_relu025*(11)+bias0_relu026*(20)+bias0_relu027*(-4)+bias0_relu028*(-8)+bias0_relu029*(44)+bias0_relu030*(-19)+bias0_relu031*(-4)+bias0_relu032*(33)+bias0_relu033*(-24)+bias0_relu034*(15)+bias0_relu035*(13)+bias0_relu036*(81)+bias0_relu037*(25)+bias0_relu038*(5)+bias0_relu039*(8)+bias0_relu040*(13)+bias0_relu041*(0)+bias0_relu042*(10)+bias0_relu043*(13)+bias0_relu044*(-58)+bias0_relu045*(-16)+bias0_relu046*(-15)+bias0_relu047*(96)+bias0_relu048*(5)+bias0_relu049*(-8)+bias0_relu050*(-4)+bias0_relu051*(21)+bias0_relu052*(21)+bias0_relu053*(-4)+bias0_relu054*(7)+bias0_relu055*(26)+bias0_relu056*(4)+bias0_relu057*(-43)+bias0_relu058*(1)+bias0_relu059*(-58)+bias0_relu060*(-26)+bias0_relu061*(20)+bias0_relu062*(-8)+bias0_relu063*(19);
assign relu0_weight27=bias0_relu00*(-62)+bias0_relu01*(60)+bias0_relu02*(-27)+bias0_relu03*(-13)+bias0_relu04*(5)+bias0_relu05*(6)+bias0_relu06*(3)+bias0_relu07*(-26)+bias0_relu08*(33)+bias0_relu09*(9)+bias0_relu010*(9)+bias0_relu011*(24)+bias0_relu012*(-13)+bias0_relu013*(-29)+bias0_relu014*(31)+bias0_relu015*(-9)+bias0_relu016*(53)+bias0_relu017*(34)+bias0_relu018*(-24)+bias0_relu019*(-17)+bias0_relu020*(20)+bias0_relu021*(-11)+bias0_relu022*(25)+bias0_relu023*(55)+bias0_relu024*(-8)+bias0_relu025*(7)+bias0_relu026*(-16)+bias0_relu027*(11)+bias0_relu028*(-6)+bias0_relu029*(-3)+bias0_relu030*(-17)+bias0_relu031*(52)+bias0_relu032*(-29)+bias0_relu033*(-13)+bias0_relu034*(27)+bias0_relu035*(44)+bias0_relu036*(-32)+bias0_relu037*(-1)+bias0_relu038*(13)+bias0_relu039*(2)+bias0_relu040*(22)+bias0_relu041*(-6)+bias0_relu042*(32)+bias0_relu043*(28)+bias0_relu044*(37)+bias0_relu045*(-19)+bias0_relu046*(39)+bias0_relu047*(10)+bias0_relu048*(36)+bias0_relu049*(-22)+bias0_relu050*(-5)+bias0_relu051*(29)+bias0_relu052*(-33)+bias0_relu053*(37)+bias0_relu054*(-16)+bias0_relu055*(0)+bias0_relu056*(25)+bias0_relu057*(-61)+bias0_relu058*(-26)+bias0_relu059*(21)+bias0_relu060*(-65)+bias0_relu061*(40)+bias0_relu062*(27)+bias0_relu063*(-7);
assign relu0_weight28=bias0_relu00*(85)+bias0_relu01*(16)+bias0_relu02*(2)+bias0_relu03*(45)+bias0_relu04*(-5)+bias0_relu05*(-2)+bias0_relu06*(-13)+bias0_relu07*(4)+bias0_relu08*(12)+bias0_relu09*(-9)+bias0_relu010*(-31)+bias0_relu011*(0)+bias0_relu012*(5)+bias0_relu013*(51)+bias0_relu014*(7)+bias0_relu015*(38)+bias0_relu016*(-3)+bias0_relu017*(-26)+bias0_relu018*(30)+bias0_relu019*(-6)+bias0_relu020*(-35)+bias0_relu021*(-17)+bias0_relu022*(11)+bias0_relu023*(5)+bias0_relu024*(-10)+bias0_relu025*(31)+bias0_relu026*(42)+bias0_relu027*(-9)+bias0_relu028*(51)+bias0_relu029*(6)+bias0_relu030*(0)+bias0_relu031*(-23)+bias0_relu032*(28)+bias0_relu033*(-2)+bias0_relu034*(-3)+bias0_relu035*(19)+bias0_relu036*(14)+bias0_relu037*(-27)+bias0_relu038*(-16)+bias0_relu039*(0)+bias0_relu040*(-20)+bias0_relu041*(35)+bias0_relu042*(0)+bias0_relu043*(-3)+bias0_relu044*(0)+bias0_relu045*(20)+bias0_relu046*(-35)+bias0_relu047*(-13)+bias0_relu048*(0)+bias0_relu049*(-3)+bias0_relu050*(24)+bias0_relu051*(12)+bias0_relu052*(76)+bias0_relu053*(2)+bias0_relu054*(-20)+bias0_relu055*(20)+bias0_relu056*(8)+bias0_relu057*(52)+bias0_relu058*(-29)+bias0_relu059*(11)+bias0_relu060*(12)+bias0_relu061*(-47)+bias0_relu062*(28)+bias0_relu063*(-9);
assign relu0_weight29=bias0_relu00*(-34)+bias0_relu01*(22)+bias0_relu02*(-12)+bias0_relu03*(25)+bias0_relu04*(17)+bias0_relu05*(6)+bias0_relu06*(15)+bias0_relu07*(-20)+bias0_relu08*(3)+bias0_relu09*(0)+bias0_relu010*(20)+bias0_relu011*(28)+bias0_relu012*(-18)+bias0_relu013*(25)+bias0_relu014*(22)+bias0_relu015*(-1)+bias0_relu016*(22)+bias0_relu017*(-25)+bias0_relu018*(20)+bias0_relu019*(-9)+bias0_relu020*(-47)+bias0_relu021*(-57)+bias0_relu022*(0)+bias0_relu023*(8)+bias0_relu024*(-25)+bias0_relu025*(15)+bias0_relu026*(43)+bias0_relu027*(10)+bias0_relu028*(-1)+bias0_relu029*(11)+bias0_relu030*(2)+bias0_relu031*(44)+bias0_relu032*(4)+bias0_relu033*(-42)+bias0_relu034*(-2)+bias0_relu035*(-3)+bias0_relu036*(3)+bias0_relu037*(-28)+bias0_relu038*(-2)+bias0_relu039*(7)+bias0_relu040*(2)+bias0_relu041*(1)+bias0_relu042*(-16)+bias0_relu043*(16)+bias0_relu044*(39)+bias0_relu045*(11)+bias0_relu046*(21)+bias0_relu047*(-2)+bias0_relu048*(26)+bias0_relu049*(13)+bias0_relu050*(-5)+bias0_relu051*(38)+bias0_relu052*(-22)+bias0_relu053*(61)+bias0_relu054*(-4)+bias0_relu055*(-3)+bias0_relu056*(26)+bias0_relu057*(-28)+bias0_relu058*(5)+bias0_relu059*(-43)+bias0_relu060*(6)+bias0_relu061*(80)+bias0_relu062*(9)+bias0_relu063*(-19);
assign relu0_weight210=bias0_relu00*(-21)+bias0_relu01*(3)+bias0_relu02*(21)+bias0_relu03*(12)+bias0_relu04*(26)+bias0_relu05*(-16)+bias0_relu06*(7)+bias0_relu07*(-21)+bias0_relu08*(27)+bias0_relu09*(-11)+bias0_relu010*(9)+bias0_relu011*(19)+bias0_relu012*(10)+bias0_relu013*(43)+bias0_relu014*(9)+bias0_relu015*(-23)+bias0_relu016*(23)+bias0_relu017*(21)+bias0_relu018*(-24)+bias0_relu019*(-5)+bias0_relu020*(-38)+bias0_relu021*(-24)+bias0_relu022*(-9)+bias0_relu023*(17)+bias0_relu024*(-33)+bias0_relu025*(27)+bias0_relu026*(56)+bias0_relu027*(-6)+bias0_relu028*(-24)+bias0_relu029*(20)+bias0_relu030*(-26)+bias0_relu031*(6)+bias0_relu032*(-28)+bias0_relu033*(-31)+bias0_relu034*(14)+bias0_relu035*(9)+bias0_relu036*(-28)+bias0_relu037*(-5)+bias0_relu038*(23)+bias0_relu039*(-6)+bias0_relu040*(19)+bias0_relu041*(8)+bias0_relu042*(46)+bias0_relu043*(-1)+bias0_relu044*(57)+bias0_relu045*(22)+bias0_relu046*(47)+bias0_relu047*(-27)+bias0_relu048*(-6)+bias0_relu049*(25)+bias0_relu050*(-24)+bias0_relu051*(-17)+bias0_relu052*(23)+bias0_relu053*(44)+bias0_relu054*(23)+bias0_relu055*(-19)+bias0_relu056*(7)+bias0_relu057*(-43)+bias0_relu058*(-31)+bias0_relu059*(-13)+bias0_relu060*(0)+bias0_relu061*(15)+bias0_relu062*(49)+bias0_relu063*(-16);
assign relu0_weight211=bias0_relu00*(14)+bias0_relu01*(-3)+bias0_relu02*(-2)+bias0_relu03*(-27)+bias0_relu04*(-26)+bias0_relu05*(0)+bias0_relu06*(0)+bias0_relu07*(19)+bias0_relu08*(-20)+bias0_relu09*(-11)+bias0_relu010*(46)+bias0_relu011*(22)+bias0_relu012*(-58)+bias0_relu013*(52)+bias0_relu014*(31)+bias0_relu015*(-18)+bias0_relu016*(49)+bias0_relu017*(20)+bias0_relu018*(-31)+bias0_relu019*(-23)+bias0_relu020*(9)+bias0_relu021*(55)+bias0_relu022*(31)+bias0_relu023*(25)+bias0_relu024*(-29)+bias0_relu025*(-8)+bias0_relu026*(60)+bias0_relu027*(10)+bias0_relu028*(-39)+bias0_relu029*(13)+bias0_relu030*(-5)+bias0_relu031*(33)+bias0_relu032*(-38)+bias0_relu033*(-8)+bias0_relu034*(9)+bias0_relu035*(-31)+bias0_relu036*(31)+bias0_relu037*(9)+bias0_relu038*(24)+bias0_relu039*(-34)+bias0_relu040*(26)+bias0_relu041*(-51)+bias0_relu042*(25)+bias0_relu043*(-16)+bias0_relu044*(11)+bias0_relu045*(42)+bias0_relu046*(-34)+bias0_relu047*(20)+bias0_relu048*(-27)+bias0_relu049*(-1)+bias0_relu050*(-11)+bias0_relu051*(-4)+bias0_relu052*(8)+bias0_relu053*(-25)+bias0_relu054*(1)+bias0_relu055*(-42)+bias0_relu056*(31)+bias0_relu057*(-25)+bias0_relu058*(-4)+bias0_relu059*(43)+bias0_relu060*(-6)+bias0_relu061*(46)+bias0_relu062*(-16)+bias0_relu063*(-26);
assign relu0_weight212=bias0_relu00*(-26)+bias0_relu01*(8)+bias0_relu02*(-13)+bias0_relu03*(29)+bias0_relu04*(-7)+bias0_relu05*(12)+bias0_relu06*(-1)+bias0_relu07*(-2)+bias0_relu08*(22)+bias0_relu09*(-7)+bias0_relu010*(0)+bias0_relu011*(-9)+bias0_relu012*(36)+bias0_relu013*(-3)+bias0_relu014*(16)+bias0_relu015*(-39)+bias0_relu016*(36)+bias0_relu017*(37)+bias0_relu018*(21)+bias0_relu019*(-3)+bias0_relu020*(-32)+bias0_relu021*(17)+bias0_relu022*(25)+bias0_relu023*(-6)+bias0_relu024*(-25)+bias0_relu025*(15)+bias0_relu026*(28)+bias0_relu027*(-12)+bias0_relu028*(-22)+bias0_relu029*(-8)+bias0_relu030*(29)+bias0_relu031*(15)+bias0_relu032*(-22)+bias0_relu033*(-14)+bias0_relu034*(-12)+bias0_relu035*(29)+bias0_relu036*(34)+bias0_relu037*(26)+bias0_relu038*(-14)+bias0_relu039*(2)+bias0_relu040*(3)+bias0_relu041*(-26)+bias0_relu042*(18)+bias0_relu043*(-10)+bias0_relu044*(-25)+bias0_relu045*(6)+bias0_relu046*(13)+bias0_relu047*(12)+bias0_relu048*(-13)+bias0_relu049*(5)+bias0_relu050*(-15)+bias0_relu051*(-16)+bias0_relu052*(26)+bias0_relu053*(-8)+bias0_relu054*(35)+bias0_relu055*(18)+bias0_relu056*(10)+bias0_relu057*(1)+bias0_relu058*(22)+bias0_relu059*(-45)+bias0_relu060*(-7)+bias0_relu061*(45)+bias0_relu062*(7)+bias0_relu063*(-25);
assign relu0_weight213=bias0_relu00*(6)+bias0_relu01*(9)+bias0_relu02*(28)+bias0_relu03*(59)+bias0_relu04*(-7)+bias0_relu05*(-8)+bias0_relu06*(7)+bias0_relu07*(0)+bias0_relu08*(-41)+bias0_relu09*(13)+bias0_relu010*(-12)+bias0_relu011*(-16)+bias0_relu012*(16)+bias0_relu013*(37)+bias0_relu014*(-6)+bias0_relu015*(-18)+bias0_relu016*(7)+bias0_relu017*(-42)+bias0_relu018*(9)+bias0_relu019*(20)+bias0_relu020*(-15)+bias0_relu021*(-40)+bias0_relu022*(-12)+bias0_relu023*(-17)+bias0_relu024*(3)+bias0_relu025*(27)+bias0_relu026*(38)+bias0_relu027*(7)+bias0_relu028*(-1)+bias0_relu029*(14)+bias0_relu030*(0)+bias0_relu031*(22)+bias0_relu032*(1)+bias0_relu033*(0)+bias0_relu034*(-20)+bias0_relu035*(10)+bias0_relu036*(21)+bias0_relu037*(-21)+bias0_relu038*(-30)+bias0_relu039*(10)+bias0_relu040*(-25)+bias0_relu041*(17)+bias0_relu042*(-19)+bias0_relu043*(-35)+bias0_relu044*(-18)+bias0_relu045*(13)+bias0_relu046*(0)+bias0_relu047*(-14)+bias0_relu048*(9)+bias0_relu049*(-6)+bias0_relu050*(0)+bias0_relu051*(9)+bias0_relu052*(-4)+bias0_relu053*(31)+bias0_relu054*(13)+bias0_relu055*(17)+bias0_relu056*(0)+bias0_relu057*(61)+bias0_relu058*(15)+bias0_relu059*(5)+bias0_relu060*(46)+bias0_relu061*(49)+bias0_relu062*(-10)+bias0_relu063*(15);
assign relu0_weight214=bias0_relu00*(8)+bias0_relu01*(-5)+bias0_relu02*(-31)+bias0_relu03*(-12)+bias0_relu04*(-11)+bias0_relu05*(31)+bias0_relu06*(-4)+bias0_relu07*(-31)+bias0_relu08*(28)+bias0_relu09*(5)+bias0_relu010*(-6)+bias0_relu011*(-8)+bias0_relu012*(1)+bias0_relu013*(-2)+bias0_relu014*(-44)+bias0_relu015*(34)+bias0_relu016*(20)+bias0_relu017*(37)+bias0_relu018*(14)+bias0_relu019*(35)+bias0_relu020*(10)+bias0_relu021*(-16)+bias0_relu022*(35)+bias0_relu023*(-6)+bias0_relu024*(-17)+bias0_relu025*(26)+bias0_relu026*(11)+bias0_relu027*(7)+bias0_relu028*(13)+bias0_relu029*(-25)+bias0_relu030*(35)+bias0_relu031*(30)+bias0_relu032*(-23)+bias0_relu033*(12)+bias0_relu034*(41)+bias0_relu035*(-31)+bias0_relu036*(-12)+bias0_relu037*(3)+bias0_relu038*(-16)+bias0_relu039*(-17)+bias0_relu040*(6)+bias0_relu041*(24)+bias0_relu042*(36)+bias0_relu043*(0)+bias0_relu044*(44)+bias0_relu045*(-63)+bias0_relu046*(9)+bias0_relu047*(-80)+bias0_relu048*(7)+bias0_relu049*(18)+bias0_relu050*(-22)+bias0_relu051*(-4)+bias0_relu052*(-7)+bias0_relu053*(-7)+bias0_relu054*(37)+bias0_relu055*(16)+bias0_relu056*(-28)+bias0_relu057*(66)+bias0_relu058*(14)+bias0_relu059*(43)+bias0_relu060*(-50)+bias0_relu061*(-2)+bias0_relu062*(-54)+bias0_relu063*(-11);
assign relu0_weight215=bias0_relu00*(15)+bias0_relu01*(25)+bias0_relu02*(32)+bias0_relu03*(-52)+bias0_relu04*(10)+bias0_relu05*(-54)+bias0_relu06*(-1)+bias0_relu07*(-7)+bias0_relu08*(-39)+bias0_relu09*(-1)+bias0_relu010*(39)+bias0_relu011*(7)+bias0_relu012*(-14)+bias0_relu013*(-12)+bias0_relu014*(-65)+bias0_relu015*(41)+bias0_relu016*(6)+bias0_relu017*(-33)+bias0_relu018*(6)+bias0_relu019*(8)+bias0_relu020*(79)+bias0_relu021*(22)+bias0_relu022*(52)+bias0_relu023*(20)+bias0_relu024*(23)+bias0_relu025*(32)+bias0_relu026*(10)+bias0_relu027*(-5)+bias0_relu028*(1)+bias0_relu029*(19)+bias0_relu030*(2)+bias0_relu031*(46)+bias0_relu032*(1)+bias0_relu033*(5)+bias0_relu034*(5)+bias0_relu035*(-7)+bias0_relu036*(39)+bias0_relu037*(9)+bias0_relu038*(-20)+bias0_relu039*(-30)+bias0_relu040*(-27)+bias0_relu041*(-9)+bias0_relu042*(-47)+bias0_relu043*(-12)+bias0_relu044*(39)+bias0_relu045*(-6)+bias0_relu046*(-4)+bias0_relu047*(1)+bias0_relu048*(4)+bias0_relu049*(-19)+bias0_relu050*(-36)+bias0_relu051*(23)+bias0_relu052*(-14)+bias0_relu053*(15)+bias0_relu054*(-9)+bias0_relu055*(22)+bias0_relu056*(-36)+bias0_relu057*(31)+bias0_relu058*(10)+bias0_relu059*(68)+bias0_relu060*(-17)+bias0_relu061*(42)+bias0_relu062*(-41)+bias0_relu063*(26);
assign relu0_weight216=bias0_relu00*(14)+bias0_relu01*(-4)+bias0_relu02*(15)+bias0_relu03*(-33)+bias0_relu04*(-19)+bias0_relu05*(12)+bias0_relu06*(-9)+bias0_relu07*(41)+bias0_relu08*(23)+bias0_relu09*(12)+bias0_relu010*(-38)+bias0_relu011*(2)+bias0_relu012*(-2)+bias0_relu013*(-25)+bias0_relu014*(-30)+bias0_relu015*(5)+bias0_relu016*(-8)+bias0_relu017*(-20)+bias0_relu018*(-25)+bias0_relu019*(2)+bias0_relu020*(-15)+bias0_relu021*(53)+bias0_relu022*(-14)+bias0_relu023*(-35)+bias0_relu024*(21)+bias0_relu025*(-21)+bias0_relu026*(-35)+bias0_relu027*(-12)+bias0_relu028*(-50)+bias0_relu029*(-38)+bias0_relu030*(21)+bias0_relu031*(12)+bias0_relu032*(-28)+bias0_relu033*(0)+bias0_relu034*(9)+bias0_relu035*(-1)+bias0_relu036*(-56)+bias0_relu037*(1)+bias0_relu038*(26)+bias0_relu039*(10)+bias0_relu040*(36)+bias0_relu041*(23)+bias0_relu042*(-33)+bias0_relu043*(-6)+bias0_relu044*(18)+bias0_relu045*(37)+bias0_relu046*(-17)+bias0_relu047*(-117)+bias0_relu048*(-16)+bias0_relu049*(38)+bias0_relu050*(6)+bias0_relu051*(15)+bias0_relu052*(0)+bias0_relu053*(7)+bias0_relu054*(33)+bias0_relu055*(3)+bias0_relu056*(31)+bias0_relu057*(42)+bias0_relu058*(37)+bias0_relu059*(26)+bias0_relu060*(14)+bias0_relu061*(-48)+bias0_relu062*(0)+bias0_relu063*(23);
assign relu0_weight217=bias0_relu00*(-23)+bias0_relu01*(34)+bias0_relu02*(5)+bias0_relu03*(-29)+bias0_relu04*(22)+bias0_relu05*(9)+bias0_relu06*(-4)+bias0_relu07*(32)+bias0_relu08*(-11)+bias0_relu09*(-1)+bias0_relu010*(-1)+bias0_relu011*(24)+bias0_relu012*(-27)+bias0_relu013*(-13)+bias0_relu014*(35)+bias0_relu015*(6)+bias0_relu016*(-48)+bias0_relu017*(-34)+bias0_relu018*(20)+bias0_relu019*(28)+bias0_relu020*(-1)+bias0_relu021*(-25)+bias0_relu022*(-5)+bias0_relu023*(32)+bias0_relu024*(29)+bias0_relu025*(12)+bias0_relu026*(-20)+bias0_relu027*(12)+bias0_relu028*(13)+bias0_relu029*(11)+bias0_relu030*(-41)+bias0_relu031*(13)+bias0_relu032*(13)+bias0_relu033*(18)+bias0_relu034*(-5)+bias0_relu035*(12)+bias0_relu036*(-7)+bias0_relu037*(-24)+bias0_relu038*(35)+bias0_relu039*(10)+bias0_relu040*(-11)+bias0_relu041*(42)+bias0_relu042*(-34)+bias0_relu043*(35)+bias0_relu044*(12)+bias0_relu045*(42)+bias0_relu046*(26)+bias0_relu047*(24)+bias0_relu048*(-14)+bias0_relu049*(42)+bias0_relu050*(30)+bias0_relu051*(-2)+bias0_relu052*(-78)+bias0_relu053*(0)+bias0_relu054*(-49)+bias0_relu055*(4)+bias0_relu056*(12)+bias0_relu057*(-54)+bias0_relu058*(-5)+bias0_relu059*(6)+bias0_relu060*(23)+bias0_relu061*(18)+bias0_relu062*(-5)+bias0_relu063*(29);
assign relu0_weight218=bias0_relu00*(14)+bias0_relu01*(11)+bias0_relu02*(-15)+bias0_relu03*(-21)+bias0_relu04*(11)+bias0_relu05*(-22)+bias0_relu06*(16)+bias0_relu07*(17)+bias0_relu08*(-76)+bias0_relu09*(-4)+bias0_relu010*(2)+bias0_relu011*(-12)+bias0_relu012*(-58)+bias0_relu013*(48)+bias0_relu014*(-24)+bias0_relu015*(15)+bias0_relu016*(-6)+bias0_relu017*(-5)+bias0_relu018*(-26)+bias0_relu019*(23)+bias0_relu020*(44)+bias0_relu021*(36)+bias0_relu022*(42)+bias0_relu023*(12)+bias0_relu024*(11)+bias0_relu025*(-11)+bias0_relu026*(-17)+bias0_relu027*(-4)+bias0_relu028*(14)+bias0_relu029*(28)+bias0_relu030*(36)+bias0_relu031*(13)+bias0_relu032*(23)+bias0_relu033*(35)+bias0_relu034*(0)+bias0_relu035*(3)+bias0_relu036*(11)+bias0_relu037*(-13)+bias0_relu038*(-11)+bias0_relu039*(-32)+bias0_relu040*(-60)+bias0_relu041*(19)+bias0_relu042*(-61)+bias0_relu043*(19)+bias0_relu044*(33)+bias0_relu045*(22)+bias0_relu046*(-13)+bias0_relu047*(27)+bias0_relu048*(16)+bias0_relu049*(15)+bias0_relu050*(8)+bias0_relu051*(22)+bias0_relu052*(-61)+bias0_relu053*(-15)+bias0_relu054*(-18)+bias0_relu055*(6)+bias0_relu056*(-5)+bias0_relu057*(-38)+bias0_relu058*(19)+bias0_relu059*(44)+bias0_relu060*(41)+bias0_relu061*(22)+bias0_relu062*(-85)+bias0_relu063*(8);
assign relu0_weight219=bias0_relu00*(72)+bias0_relu01*(-21)+bias0_relu02*(15)+bias0_relu03*(59)+bias0_relu04*(-10)+bias0_relu05*(25)+bias0_relu06*(-3)+bias0_relu07*(3)+bias0_relu08*(7)+bias0_relu09*(5)+bias0_relu010*(-14)+bias0_relu011*(-17)+bias0_relu012*(-16)+bias0_relu013*(15)+bias0_relu014*(24)+bias0_relu015*(22)+bias0_relu016*(-14)+bias0_relu017*(23)+bias0_relu018*(23)+bias0_relu019*(8)+bias0_relu020*(-11)+bias0_relu021*(44)+bias0_relu022*(-40)+bias0_relu023*(-26)+bias0_relu024*(-4)+bias0_relu025*(-34)+bias0_relu026*(18)+bias0_relu027*(13)+bias0_relu028*(0)+bias0_relu029*(-3)+bias0_relu030*(46)+bias0_relu031*(-18)+bias0_relu032*(-29)+bias0_relu033*(22)+bias0_relu034*(-16)+bias0_relu035*(26)+bias0_relu036*(30)+bias0_relu037*(13)+bias0_relu038*(-15)+bias0_relu039*(0)+bias0_relu040*(0)+bias0_relu041*(-53)+bias0_relu042*(-1)+bias0_relu043*(-8)+bias0_relu044*(-33)+bias0_relu045*(-14)+bias0_relu046*(-73)+bias0_relu047*(1)+bias0_relu048*(-13)+bias0_relu049*(-9)+bias0_relu050*(33)+bias0_relu051*(-2)+bias0_relu052*(60)+bias0_relu053*(-32)+bias0_relu054*(24)+bias0_relu055*(14)+bias0_relu056*(20)+bias0_relu057*(37)+bias0_relu058*(36)+bias0_relu059*(-16)+bias0_relu060*(37)+bias0_relu061*(23)+bias0_relu062*(4)+bias0_relu063*(3);
assign relu0_weight220=bias0_relu00*(-15)+bias0_relu01*(-53)+bias0_relu02*(-19)+bias0_relu03*(-36)+bias0_relu04*(-18)+bias0_relu05*(-11)+bias0_relu06*(11)+bias0_relu07*(21)+bias0_relu08*(6)+bias0_relu09*(16)+bias0_relu010*(20)+bias0_relu011*(-16)+bias0_relu012*(18)+bias0_relu013*(-20)+bias0_relu014*(-36)+bias0_relu015*(31)+bias0_relu016*(9)+bias0_relu017*(24)+bias0_relu018*(-9)+bias0_relu019*(48)+bias0_relu020*(39)+bias0_relu021*(29)+bias0_relu022*(1)+bias0_relu023*(-24)+bias0_relu024*(-6)+bias0_relu025*(22)+bias0_relu026*(-8)+bias0_relu027*(10)+bias0_relu028*(29)+bias0_relu029*(-25)+bias0_relu030*(17)+bias0_relu031*(25)+bias0_relu032*(19)+bias0_relu033*(15)+bias0_relu034*(27)+bias0_relu035*(-10)+bias0_relu036*(12)+bias0_relu037*(22)+bias0_relu038*(-20)+bias0_relu039*(16)+bias0_relu040*(8)+bias0_relu041*(14)+bias0_relu042*(7)+bias0_relu043*(-34)+bias0_relu044*(10)+bias0_relu045*(-25)+bias0_relu046*(4)+bias0_relu047*(-48)+bias0_relu048*(21)+bias0_relu049*(2)+bias0_relu050*(0)+bias0_relu051*(7)+bias0_relu052*(-58)+bias0_relu053*(5)+bias0_relu054*(15)+bias0_relu055*(20)+bias0_relu056*(-1)+bias0_relu057*(68)+bias0_relu058*(20)+bias0_relu059*(53)+bias0_relu060*(11)+bias0_relu061*(1)+bias0_relu062*(-36)+bias0_relu063*(4);
assign relu0_weight221=bias0_relu00*(-9)+bias0_relu01*(4)+bias0_relu02*(42)+bias0_relu03*(4)+bias0_relu04*(7)+bias0_relu05*(-26)+bias0_relu06*(-10)+bias0_relu07*(-16)+bias0_relu08*(30)+bias0_relu09*(11)+bias0_relu010*(0)+bias0_relu011*(9)+bias0_relu012*(9)+bias0_relu013*(46)+bias0_relu014*(7)+bias0_relu015*(-39)+bias0_relu016*(47)+bias0_relu017*(53)+bias0_relu018*(-64)+bias0_relu019*(-5)+bias0_relu020*(41)+bias0_relu021*(26)+bias0_relu022*(25)+bias0_relu023*(-3)+bias0_relu024*(-3)+bias0_relu025*(-19)+bias0_relu026*(35)+bias0_relu027*(-3)+bias0_relu028*(-34)+bias0_relu029*(4)+bias0_relu030*(8)+bias0_relu031*(36)+bias0_relu032*(-11)+bias0_relu033*(25)+bias0_relu034*(-17)+bias0_relu035*(9)+bias0_relu036*(-50)+bias0_relu037*(0)+bias0_relu038*(-13)+bias0_relu039*(-17)+bias0_relu040*(13)+bias0_relu041*(5)+bias0_relu042*(29)+bias0_relu043*(-9)+bias0_relu044*(73)+bias0_relu045*(14)+bias0_relu046*(39)+bias0_relu047*(-54)+bias0_relu048*(14)+bias0_relu049*(7)+bias0_relu050*(-14)+bias0_relu051*(-29)+bias0_relu052*(20)+bias0_relu053*(4)+bias0_relu054*(15)+bias0_relu055*(-7)+bias0_relu056*(-25)+bias0_relu057*(16)+bias0_relu058*(-37)+bias0_relu059*(27)+bias0_relu060*(-1)+bias0_relu061*(14)+bias0_relu062*(8)+bias0_relu063*(-18);
assign relu0_weight222=bias0_relu00*(32)+bias0_relu01*(-10)+bias0_relu02*(-18)+bias0_relu03*(17)+bias0_relu04*(28)+bias0_relu05*(-8)+bias0_relu06*(-1)+bias0_relu07*(28)+bias0_relu08*(-5)+bias0_relu09*(15)+bias0_relu010*(9)+bias0_relu011*(-5)+bias0_relu012*(33)+bias0_relu013*(21)+bias0_relu014*(22)+bias0_relu015*(-40)+bias0_relu016*(59)+bias0_relu017*(27)+bias0_relu018*(7)+bias0_relu019*(-3)+bias0_relu020*(45)+bias0_relu021*(35)+bias0_relu022*(-23)+bias0_relu023*(23)+bias0_relu024*(20)+bias0_relu025*(25)+bias0_relu026*(28)+bias0_relu027*(-9)+bias0_relu028*(-19)+bias0_relu029*(22)+bias0_relu030*(10)+bias0_relu031*(-18)+bias0_relu032*(30)+bias0_relu033*(44)+bias0_relu034*(1)+bias0_relu035*(-33)+bias0_relu036*(7)+bias0_relu037*(56)+bias0_relu038*(-6)+bias0_relu039*(-20)+bias0_relu040*(5)+bias0_relu041*(-9)+bias0_relu042*(43)+bias0_relu043*(-7)+bias0_relu044*(-25)+bias0_relu045*(15)+bias0_relu046*(15)+bias0_relu047*(83)+bias0_relu048*(-11)+bias0_relu049*(13)+bias0_relu050*(4)+bias0_relu051*(-25)+bias0_relu052*(42)+bias0_relu053*(-35)+bias0_relu054*(27)+bias0_relu055*(18)+bias0_relu056*(0)+bias0_relu057*(-18)+bias0_relu058*(-34)+bias0_relu059*(-14)+bias0_relu060*(31)+bias0_relu061*(-6)+bias0_relu062*(-8)+bias0_relu063*(-15);
assign relu0_weight223=bias0_relu00*(-43)+bias0_relu01*(-12)+bias0_relu02*(8)+bias0_relu03*(12)+bias0_relu04*(31)+bias0_relu05*(0)+bias0_relu06*(14)+bias0_relu07*(-8)+bias0_relu08*(6)+bias0_relu09*(-14)+bias0_relu010*(38)+bias0_relu011*(-10)+bias0_relu012*(-3)+bias0_relu013*(3)+bias0_relu014*(-4)+bias0_relu015*(-30)+bias0_relu016*(23)+bias0_relu017*(-21)+bias0_relu018*(0)+bias0_relu019*(18)+bias0_relu020*(-20)+bias0_relu021*(-37)+bias0_relu022*(11)+bias0_relu023*(14)+bias0_relu024*(-3)+bias0_relu025*(27)+bias0_relu026*(39)+bias0_relu027*(-5)+bias0_relu028*(-7)+bias0_relu029*(36)+bias0_relu030*(19)+bias0_relu031*(23)+bias0_relu032*(30)+bias0_relu033*(-39)+bias0_relu034*(-21)+bias0_relu035*(0)+bias0_relu036*(37)+bias0_relu037*(-6)+bias0_relu038*(2)+bias0_relu039*(-12)+bias0_relu040*(-5)+bias0_relu041*(-13)+bias0_relu042*(-9)+bias0_relu043*(-22)+bias0_relu044*(3)+bias0_relu045*(-21)+bias0_relu046*(34)+bias0_relu047*(8)+bias0_relu048*(9)+bias0_relu049*(-2)+bias0_relu050*(3)+bias0_relu051*(34)+bias0_relu052*(-49)+bias0_relu053*(50)+bias0_relu054*(13)+bias0_relu055*(21)+bias0_relu056*(9)+bias0_relu057*(12)+bias0_relu058*(22)+bias0_relu059*(-25)+bias0_relu060*(0)+bias0_relu061*(73)+bias0_relu062*(1)+bias0_relu063*(14);
assign relu0_weight224=bias0_relu00*(16)+bias0_relu01*(18)+bias0_relu02*(-28)+bias0_relu03*(-18)+bias0_relu04*(25)+bias0_relu05*(-16)+bias0_relu06*(16)+bias0_relu07*(-20)+bias0_relu08*(34)+bias0_relu09*(-10)+bias0_relu010*(20)+bias0_relu011*(-9)+bias0_relu012*(-4)+bias0_relu013*(-11)+bias0_relu014*(-25)+bias0_relu015*(41)+bias0_relu016*(32)+bias0_relu017*(7)+bias0_relu018*(7)+bias0_relu019*(0)+bias0_relu020*(31)+bias0_relu021*(17)+bias0_relu022*(53)+bias0_relu023*(18)+bias0_relu024*(-19)+bias0_relu025*(41)+bias0_relu026*(-21)+bias0_relu027*(-1)+bias0_relu028*(32)+bias0_relu029*(3)+bias0_relu030*(8)+bias0_relu031*(25)+bias0_relu032*(-19)+bias0_relu033*(36)+bias0_relu034*(55)+bias0_relu035*(37)+bias0_relu036*(26)+bias0_relu037*(48)+bias0_relu038*(-6)+bias0_relu039*(8)+bias0_relu040*(17)+bias0_relu041*(22)+bias0_relu042*(40)+bias0_relu043*(1)+bias0_relu044*(9)+bias0_relu045*(-39)+bias0_relu046*(-12)+bias0_relu047*(27)+bias0_relu048*(34)+bias0_relu049*(-33)+bias0_relu050*(-15)+bias0_relu051*(2)+bias0_relu052*(33)+bias0_relu053*(-3)+bias0_relu054*(-3)+bias0_relu055*(10)+bias0_relu056*(4)+bias0_relu057*(-2)+bias0_relu058*(-9)+bias0_relu059*(34)+bias0_relu060*(-23)+bias0_relu061*(34)+bias0_relu062*(-6)+bias0_relu063*(-7);
assign relu0_weight225=bias0_relu00*(21)+bias0_relu01*(25)+bias0_relu02*(49)+bias0_relu03*(-11)+bias0_relu04*(-4)+bias0_relu05*(-26)+bias0_relu06*(15)+bias0_relu07*(13)+bias0_relu08*(-5)+bias0_relu09*(-9)+bias0_relu010*(-6)+bias0_relu011*(-5)+bias0_relu012*(-4)+bias0_relu013*(55)+bias0_relu014*(-16)+bias0_relu015*(-56)+bias0_relu016*(18)+bias0_relu017*(23)+bias0_relu018*(-55)+bias0_relu019*(56)+bias0_relu020*(33)+bias0_relu021*(28)+bias0_relu022*(-12)+bias0_relu023*(-29)+bias0_relu024*(22)+bias0_relu025*(-13)+bias0_relu026*(-11)+bias0_relu027*(-4)+bias0_relu028*(-16)+bias0_relu029*(-6)+bias0_relu030*(13)+bias0_relu031*(31)+bias0_relu032*(-11)+bias0_relu033*(31)+bias0_relu034*(-27)+bias0_relu035*(26)+bias0_relu036*(-67)+bias0_relu037*(-11)+bias0_relu038*(16)+bias0_relu039*(6)+bias0_relu040*(5)+bias0_relu041*(35)+bias0_relu042*(-23)+bias0_relu043*(-8)+bias0_relu044*(26)+bias0_relu045*(23)+bias0_relu046*(7)+bias0_relu047*(-23)+bias0_relu048*(9)+bias0_relu049*(15)+bias0_relu050*(9)+bias0_relu051*(4)+bias0_relu052*(-11)+bias0_relu053*(48)+bias0_relu054*(13)+bias0_relu055*(-10)+bias0_relu056*(10)+bias0_relu057*(19)+bias0_relu058*(4)+bias0_relu059*(72)+bias0_relu060*(3)+bias0_relu061*(1)+bias0_relu062*(0)+bias0_relu063*(18);
assign relu0_weight226=bias0_relu00*(12)+bias0_relu01*(1)+bias0_relu02*(1)+bias0_relu03*(-6)+bias0_relu04*(0)+bias0_relu05*(-14)+bias0_relu06*(8)+bias0_relu07*(-6)+bias0_relu08*(-16)+bias0_relu09*(-5)+bias0_relu010*(-7)+bias0_relu011*(-11)+bias0_relu012*(-5)+bias0_relu013*(-13)+bias0_relu014*(-4)+bias0_relu015*(6)+bias0_relu016*(2)+bias0_relu017*(-3)+bias0_relu018*(-10)+bias0_relu019*(-16)+bias0_relu020*(0)+bias0_relu021*(-14)+bias0_relu022*(-4)+bias0_relu023*(-6)+bias0_relu024*(3)+bias0_relu025*(-14)+bias0_relu026*(-14)+bias0_relu027*(12)+bias0_relu028*(-10)+bias0_relu029*(-11)+bias0_relu030*(-12)+bias0_relu031*(-8)+bias0_relu032*(-12)+bias0_relu033*(-6)+bias0_relu034*(2)+bias0_relu035*(-9)+bias0_relu036*(5)+bias0_relu037*(3)+bias0_relu038*(2)+bias0_relu039*(6)+bias0_relu040*(-1)+bias0_relu041*(-4)+bias0_relu042*(-9)+bias0_relu043*(7)+bias0_relu044*(14)+bias0_relu045*(-18)+bias0_relu046*(3)+bias0_relu047*(-1)+bias0_relu048*(11)+bias0_relu049*(-18)+bias0_relu050*(11)+bias0_relu051*(-2)+bias0_relu052*(-3)+bias0_relu053*(4)+bias0_relu054*(-2)+bias0_relu055*(-9)+bias0_relu056*(-12)+bias0_relu057*(-8)+bias0_relu058*(9)+bias0_relu059*(-7)+bias0_relu060*(-9)+bias0_relu061*(-5)+bias0_relu062*(-11)+bias0_relu063*(-7);
assign relu0_weight227=bias0_relu00*(-45)+bias0_relu01*(-14)+bias0_relu02*(-59)+bias0_relu03*(-15)+bias0_relu04*(-5)+bias0_relu05*(-3)+bias0_relu06*(5)+bias0_relu07*(28)+bias0_relu08*(-10)+bias0_relu09*(2)+bias0_relu010*(24)+bias0_relu011*(7)+bias0_relu012*(19)+bias0_relu013*(-28)+bias0_relu014*(1)+bias0_relu015*(16)+bias0_relu016*(-31)+bias0_relu017*(-9)+bias0_relu018*(29)+bias0_relu019*(7)+bias0_relu020*(1)+bias0_relu021*(-5)+bias0_relu022*(26)+bias0_relu023*(6)+bias0_relu024*(7)+bias0_relu025*(-4)+bias0_relu026*(-34)+bias0_relu027*(5)+bias0_relu028*(6)+bias0_relu029*(27)+bias0_relu030*(19)+bias0_relu031*(6)+bias0_relu032*(18)+bias0_relu033*(19)+bias0_relu034*(29)+bias0_relu035*(-22)+bias0_relu036*(79)+bias0_relu037*(42)+bias0_relu038*(6)+bias0_relu039*(8)+bias0_relu040*(20)+bias0_relu041*(-13)+bias0_relu042*(0)+bias0_relu043*(5)+bias0_relu044*(-67)+bias0_relu045*(25)+bias0_relu046*(-31)+bias0_relu047*(90)+bias0_relu048*(-4)+bias0_relu049*(20)+bias0_relu050*(0)+bias0_relu051*(11)+bias0_relu052*(-41)+bias0_relu053*(-54)+bias0_relu054*(8)+bias0_relu055*(6)+bias0_relu056*(22)+bias0_relu057*(-10)+bias0_relu058*(-19)+bias0_relu059*(-8)+bias0_relu060*(37)+bias0_relu061*(5)+bias0_relu062*(9)+bias0_relu063*(27);
assign relu0_weight228=bias0_relu00*(12)+bias0_relu01*(10)+bias0_relu02*(39)+bias0_relu03*(-33)+bias0_relu04*(21)+bias0_relu05*(-3)+bias0_relu06*(7)+bias0_relu07*(17)+bias0_relu08*(-9)+bias0_relu09*(-11)+bias0_relu010*(-5)+bias0_relu011*(19)+bias0_relu012*(-42)+bias0_relu013*(12)+bias0_relu014*(-3)+bias0_relu015*(38)+bias0_relu016*(-35)+bias0_relu017*(-57)+bias0_relu018*(3)+bias0_relu019*(17)+bias0_relu020*(11)+bias0_relu021*(-54)+bias0_relu022*(12)+bias0_relu023*(22)+bias0_relu024*(-3)+bias0_relu025*(13)+bias0_relu026*(-22)+bias0_relu027*(-6)+bias0_relu028*(33)+bias0_relu029*(14)+bias0_relu030*(-32)+bias0_relu031*(6)+bias0_relu032*(29)+bias0_relu033*(-10)+bias0_relu034*(-22)+bias0_relu035*(22)+bias0_relu036*(-8)+bias0_relu037*(-47)+bias0_relu038*(5)+bias0_relu039*(10)+bias0_relu040*(-7)+bias0_relu041*(52)+bias0_relu042*(-41)+bias0_relu043*(30)+bias0_relu044*(41)+bias0_relu045*(28)+bias0_relu046*(14)+bias0_relu047*(0)+bias0_relu048*(15)+bias0_relu049*(20)+bias0_relu050*(13)+bias0_relu051*(18)+bias0_relu052*(-52)+bias0_relu053*(33)+bias0_relu054*(-40)+bias0_relu055*(-2)+bias0_relu056*(18)+bias0_relu057*(-11)+bias0_relu058*(1)+bias0_relu059*(10)+bias0_relu060*(-10)+bias0_relu061*(-1)+bias0_relu062*(-20)+bias0_relu063*(26);
assign relu0_weight229=bias0_relu00*(40)+bias0_relu01*(-29)+bias0_relu02*(29)+bias0_relu03*(30)+bias0_relu04*(-2)+bias0_relu05*(28)+bias0_relu06*(4)+bias0_relu07*(-11)+bias0_relu08*(8)+bias0_relu09*(-8)+bias0_relu010*(5)+bias0_relu011*(18)+bias0_relu012*(-21)+bias0_relu013*(23)+bias0_relu014*(12)+bias0_relu015*(40)+bias0_relu016*(-43)+bias0_relu017*(-32)+bias0_relu018*(21)+bias0_relu019*(-1)+bias0_relu020*(-55)+bias0_relu021*(-48)+bias0_relu022*(-20)+bias0_relu023*(-8)+bias0_relu024*(4)+bias0_relu025*(-2)+bias0_relu026*(36)+bias0_relu027*(6)+bias0_relu028*(32)+bias0_relu029*(18)+bias0_relu030*(-27)+bias0_relu031*(-65)+bias0_relu032*(29)+bias0_relu033*(-11)+bias0_relu034*(31)+bias0_relu035*(12)+bias0_relu036*(6)+bias0_relu037*(-45)+bias0_relu038*(-4)+bias0_relu039*(12)+bias0_relu040*(-1)+bias0_relu041*(27)+bias0_relu042*(-9)+bias0_relu043*(29)+bias0_relu044*(29)+bias0_relu045*(9)+bias0_relu046*(-4)+bias0_relu047*(-14)+bias0_relu048*(23)+bias0_relu049*(-6)+bias0_relu050*(28)+bias0_relu051*(-3)+bias0_relu052*(44)+bias0_relu053*(18)+bias0_relu054*(-18)+bias0_relu055*(4)+bias0_relu056*(20)+bias0_relu057*(13)+bias0_relu058*(0)+bias0_relu059*(-27)+bias0_relu060*(24)+bias0_relu061*(-68)+bias0_relu062*(18)+bias0_relu063*(11);
assign relu0_weight230=bias0_relu00*(99)+bias0_relu01*(21)+bias0_relu02*(8)+bias0_relu03*(10)+bias0_relu04*(0)+bias0_relu05*(22)+bias0_relu06*(3)+bias0_relu07*(21)+bias0_relu08*(40)+bias0_relu09*(12)+bias0_relu010*(-17)+bias0_relu011*(15)+bias0_relu012*(-15)+bias0_relu013*(14)+bias0_relu014*(12)+bias0_relu015*(40)+bias0_relu016*(17)+bias0_relu017*(-13)+bias0_relu018*(25)+bias0_relu019*(-23)+bias0_relu020*(7)+bias0_relu021*(-15)+bias0_relu022*(5)+bias0_relu023*(4)+bias0_relu024*(14)+bias0_relu025*(-1)+bias0_relu026*(-12)+bias0_relu027*(6)+bias0_relu028*(25)+bias0_relu029*(15)+bias0_relu030*(-32)+bias0_relu031*(-20)+bias0_relu032*(-3)+bias0_relu033*(-6)+bias0_relu034*(-12)+bias0_relu035*(36)+bias0_relu036*(-6)+bias0_relu037*(-16)+bias0_relu038*(-2)+bias0_relu039*(-9)+bias0_relu040*(35)+bias0_relu041*(15)+bias0_relu042*(-3)+bias0_relu043*(2)+bias0_relu044*(19)+bias0_relu045*(-1)+bias0_relu046*(-20)+bias0_relu047*(24)+bias0_relu048*(9)+bias0_relu049*(-12)+bias0_relu050*(-11)+bias0_relu051*(7)+bias0_relu052*(82)+bias0_relu053*(-10)+bias0_relu054*(17)+bias0_relu055*(-5)+bias0_relu056*(17)+bias0_relu057*(14)+bias0_relu058*(-4)+bias0_relu059*(-5)+bias0_relu060*(-54)+bias0_relu061*(-39)+bias0_relu062*(6)+bias0_relu063*(19);
assign relu0_weight231=bias0_relu00*(0)+bias0_relu01*(-14)+bias0_relu02*(-24)+bias0_relu03*(-2)+bias0_relu04*(-23)+bias0_relu05*(19)+bias0_relu06*(-6)+bias0_relu07*(16)+bias0_relu08*(6)+bias0_relu09*(-9)+bias0_relu010*(8)+bias0_relu011*(-1)+bias0_relu012*(15)+bias0_relu013*(-19)+bias0_relu014*(-15)+bias0_relu015*(36)+bias0_relu016*(-32)+bias0_relu017*(-27)+bias0_relu018*(58)+bias0_relu019*(-19)+bias0_relu020*(-7)+bias0_relu021*(38)+bias0_relu022*(34)+bias0_relu023*(0)+bias0_relu024*(15)+bias0_relu025*(2)+bias0_relu026*(-32)+bias0_relu027*(15)+bias0_relu028*(-12)+bias0_relu029*(3)+bias0_relu030*(15)+bias0_relu031*(-15)+bias0_relu032*(-7)+bias0_relu033*(15)+bias0_relu034*(27)+bias0_relu035*(16)+bias0_relu036*(65)+bias0_relu037*(31)+bias0_relu038*(12)+bias0_relu039*(8)+bias0_relu040*(23)+bias0_relu041*(-6)+bias0_relu042*(-6)+bias0_relu043*(7)+bias0_relu044*(-56)+bias0_relu045*(-17)+bias0_relu046*(-44)+bias0_relu047*(42)+bias0_relu048*(3)+bias0_relu049*(0)+bias0_relu050*(8)+bias0_relu051*(-16)+bias0_relu052*(27)+bias0_relu053*(-52)+bias0_relu054*(16)+bias0_relu055*(-15)+bias0_relu056*(26)+bias0_relu057*(27)+bias0_relu058*(12)+bias0_relu059*(10)+bias0_relu060*(18)+bias0_relu061*(-12)+bias0_relu062*(12)+bias0_relu063*(24);
wire [DATAWIDTH-1:0]   weight2_bias20;
wire [DATAWIDTH-1:0]   weight2_bias21;
wire [DATAWIDTH-1:0]   weight2_bias22;
wire [DATAWIDTH-1:0]   weight2_bias23;
wire [DATAWIDTH-1:0]   weight2_bias24;
wire [DATAWIDTH-1:0]   weight2_bias25;
wire [DATAWIDTH-1:0]   weight2_bias26;
wire [DATAWIDTH-1:0]   weight2_bias27;
wire [DATAWIDTH-1:0]   weight2_bias28;
wire [DATAWIDTH-1:0]   weight2_bias29;
wire [DATAWIDTH-1:0]   weight2_bias210;
wire [DATAWIDTH-1:0]   weight2_bias211;
wire [DATAWIDTH-1:0]   weight2_bias212;
wire [DATAWIDTH-1:0]   weight2_bias213;
wire [DATAWIDTH-1:0]   weight2_bias214;
wire [DATAWIDTH-1:0]   weight2_bias215;
wire [DATAWIDTH-1:0]   weight2_bias216;
wire [DATAWIDTH-1:0]   weight2_bias217;
wire [DATAWIDTH-1:0]   weight2_bias218;
wire [DATAWIDTH-1:0]   weight2_bias219;
wire [DATAWIDTH-1:0]   weight2_bias220;
wire [DATAWIDTH-1:0]   weight2_bias221;
wire [DATAWIDTH-1:0]   weight2_bias222;
wire [DATAWIDTH-1:0]   weight2_bias223;
wire [DATAWIDTH-1:0]   weight2_bias224;
wire [DATAWIDTH-1:0]   weight2_bias225;
wire [DATAWIDTH-1:0]   weight2_bias226;
wire [DATAWIDTH-1:0]   weight2_bias227;
wire [DATAWIDTH-1:0]   weight2_bias228;
wire [DATAWIDTH-1:0]   weight2_bias229;
wire [DATAWIDTH-1:0]   weight2_bias230;
wire [DATAWIDTH-1:0]   weight2_bias231;
assign weight2_bias20=relu0_weight20+(-28);
assign weight2_bias21=relu0_weight21+(27);
assign weight2_bias22=relu0_weight22+(9);
assign weight2_bias23=relu0_weight23+(7);
assign weight2_bias24=relu0_weight24+(3);
assign weight2_bias25=relu0_weight25+(24);
assign weight2_bias26=relu0_weight26+(7);
assign weight2_bias27=relu0_weight27+(0);
assign weight2_bias28=relu0_weight28+(31);
assign weight2_bias29=relu0_weight29+(-21);
assign weight2_bias210=relu0_weight210+(-15);
assign weight2_bias211=relu0_weight211+(-20);
assign weight2_bias212=relu0_weight212+(-14);
assign weight2_bias213=relu0_weight213+(-13);
assign weight2_bias214=relu0_weight214+(13);
assign weight2_bias215=relu0_weight215+(4);
assign weight2_bias216=relu0_weight216+(12);
assign weight2_bias217=relu0_weight217+(30);
assign weight2_bias218=relu0_weight218+(6);
assign weight2_bias219=relu0_weight219+(-9);
assign weight2_bias220=relu0_weight220+(12);
assign weight2_bias221=relu0_weight221+(24);
assign weight2_bias222=relu0_weight222+(30);
assign weight2_bias223=relu0_weight223+(-9);
assign weight2_bias224=relu0_weight224+(34);
assign weight2_bias225=relu0_weight225+(16);
assign weight2_bias226=relu0_weight226+(-17);
assign weight2_bias227=relu0_weight227+(10);
assign weight2_bias228=relu0_weight228+(3);
assign weight2_bias229=relu0_weight229+(38);
assign weight2_bias230=relu0_weight230+(7);
assign weight2_bias231=relu0_weight231+(19);
wire [DATAWIDTH-1:0]   bias2_relu20;
wire [DATAWIDTH-1:0]   bias2_relu21;
wire [DATAWIDTH-1:0]   bias2_relu22;
wire [DATAWIDTH-1:0]   bias2_relu23;
wire [DATAWIDTH-1:0]   bias2_relu24;
wire [DATAWIDTH-1:0]   bias2_relu25;
wire [DATAWIDTH-1:0]   bias2_relu26;
wire [DATAWIDTH-1:0]   bias2_relu27;
wire [DATAWIDTH-1:0]   bias2_relu28;
wire [DATAWIDTH-1:0]   bias2_relu29;
wire [DATAWIDTH-1:0]   bias2_relu210;
wire [DATAWIDTH-1:0]   bias2_relu211;
wire [DATAWIDTH-1:0]   bias2_relu212;
wire [DATAWIDTH-1:0]   bias2_relu213;
wire [DATAWIDTH-1:0]   bias2_relu214;
wire [DATAWIDTH-1:0]   bias2_relu215;
wire [DATAWIDTH-1:0]   bias2_relu216;
wire [DATAWIDTH-1:0]   bias2_relu217;
wire [DATAWIDTH-1:0]   bias2_relu218;
wire [DATAWIDTH-1:0]   bias2_relu219;
wire [DATAWIDTH-1:0]   bias2_relu220;
wire [DATAWIDTH-1:0]   bias2_relu221;
wire [DATAWIDTH-1:0]   bias2_relu222;
wire [DATAWIDTH-1:0]   bias2_relu223;
wire [DATAWIDTH-1:0]   bias2_relu224;
wire [DATAWIDTH-1:0]   bias2_relu225;
wire [DATAWIDTH-1:0]   bias2_relu226;
wire [DATAWIDTH-1:0]   bias2_relu227;
wire [DATAWIDTH-1:0]   bias2_relu228;
wire [DATAWIDTH-1:0]   bias2_relu229;
wire [DATAWIDTH-1:0]   bias2_relu230;
wire [DATAWIDTH-1:0]   bias2_relu231;
assign bias2_relu20=(weight2_bias20[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias20;
assign bias2_relu21=(weight2_bias21[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias21;
assign bias2_relu22=(weight2_bias22[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias22;
assign bias2_relu23=(weight2_bias23[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias23;
assign bias2_relu24=(weight2_bias24[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias24;
assign bias2_relu25=(weight2_bias25[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias25;
assign bias2_relu26=(weight2_bias26[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias26;
assign bias2_relu27=(weight2_bias27[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias27;
assign bias2_relu28=(weight2_bias28[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias28;
assign bias2_relu29=(weight2_bias29[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias29;
assign bias2_relu210=(weight2_bias210[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias210;
assign bias2_relu211=(weight2_bias211[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias211;
assign bias2_relu212=(weight2_bias212[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias212;
assign bias2_relu213=(weight2_bias213[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias213;
assign bias2_relu214=(weight2_bias214[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias214;
assign bias2_relu215=(weight2_bias215[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias215;
assign bias2_relu216=(weight2_bias216[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias216;
assign bias2_relu217=(weight2_bias217[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias217;
assign bias2_relu218=(weight2_bias218[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias218;
assign bias2_relu219=(weight2_bias219[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias219;
assign bias2_relu220=(weight2_bias220[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias220;
assign bias2_relu221=(weight2_bias221[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias221;
assign bias2_relu222=(weight2_bias222[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias222;
assign bias2_relu223=(weight2_bias223[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias223;
assign bias2_relu224=(weight2_bias224[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias224;
assign bias2_relu225=(weight2_bias225[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias225;
assign bias2_relu226=(weight2_bias226[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias226;
assign bias2_relu227=(weight2_bias227[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias227;
assign bias2_relu228=(weight2_bias228[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias228;
assign bias2_relu229=(weight2_bias229[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias229;
assign bias2_relu230=(weight2_bias230[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias230;
assign bias2_relu231=(weight2_bias231[DATAWIDTH-1]==1'b1)   ?   {DATAWIDTH{1'b0}}:weight2_bias231;

wire [DATAWIDTH-1:0]   relu2_weight40;
wire [DATAWIDTH-1:0]   relu2_weight41;
wire [DATAWIDTH-1:0]   relu2_weight42;
wire [DATAWIDTH-1:0]   relu2_weight43;
wire [DATAWIDTH-1:0]   relu2_weight44;
wire [DATAWIDTH-1:0]   relu2_weight45;
wire [DATAWIDTH-1:0]   relu2_weight46;
wire [DATAWIDTH-1:0]   relu2_weight47;
wire [DATAWIDTH-1:0]   relu2_weight48;
wire [DATAWIDTH-1:0]   relu2_weight49;
assign relu2_weight40=bias2_relu20*(29)+bias2_relu21*(27)+bias2_relu22*(12)+bias2_relu23*(14)+bias2_relu24*(32)+bias2_relu25*(0)+bias2_relu26*(-71)+bias2_relu27*(-7)+bias2_relu28*(-49)+bias2_relu29*(1)+bias2_relu210*(-45)+bias2_relu211*(-80)+bias2_relu212*(11)+bias2_relu213*(-19)+bias2_relu214*(17)+bias2_relu215*(-44)+bias2_relu216*(45)+bias2_relu217*(-27)+bias2_relu218*(-6)+bias2_relu219*(29)+bias2_relu220*(16)+bias2_relu221*(10)+bias2_relu222*(-55)+bias2_relu223*(-56)+bias2_relu224*(0)+bias2_relu225*(19)+bias2_relu226*(-3)+bias2_relu227*(-3)+bias2_relu228*(-15)+bias2_relu229*(-30)+bias2_relu230*(-36)+bias2_relu231*(31);
assign relu2_weight41=bias2_relu20*(-30)+bias2_relu21*(-50)+bias2_relu22*(-48)+bias2_relu23*(-79)+bias2_relu24*(-24)+bias2_relu25*(-93)+bias2_relu26*(10)+bias2_relu27*(49)+bias2_relu28*(46)+bias2_relu29*(41)+bias2_relu210*(33)+bias2_relu211*(43)+bias2_relu212*(23)+bias2_relu213*(-1)+bias2_relu214*(52)+bias2_relu215*(26)+bias2_relu216*(25)+bias2_relu217*(-28)+bias2_relu218*(-50)+bias2_relu219*(-13)+bias2_relu220*(-41)+bias2_relu221*(14)+bias2_relu222*(-23)+bias2_relu223*(9)+bias2_relu224*(24)+bias2_relu225*(-53)+bias2_relu226*(12)+bias2_relu227*(-36)+bias2_relu228*(10)+bias2_relu229*(24)+bias2_relu230*(39)+bias2_relu231*(-31);
assign relu2_weight42=bias2_relu20*(-1)+bias2_relu21*(34)+bias2_relu22*(24)+bias2_relu23*(-26)+bias2_relu24*(30)+bias2_relu25*(-19)+bias2_relu26*(-46)+bias2_relu27*(34)+bias2_relu28*(-44)+bias2_relu29*(-2)+bias2_relu210*(34)+bias2_relu211*(34)+bias2_relu212*(0)+bias2_relu213*(-20)+bias2_relu214*(-57)+bias2_relu215*(-5)+bias2_relu216*(-47)+bias2_relu217*(18)+bias2_relu218*(37)+bias2_relu219*(-22)+bias2_relu220*(-24)+bias2_relu221*(63)+bias2_relu222*(30)+bias2_relu223*(-14)+bias2_relu224*(-18)+bias2_relu225*(41)+bias2_relu226*(-3)+bias2_relu227*(-9)+bias2_relu228*(-6)+bias2_relu229*(-41)+bias2_relu230*(-26)+bias2_relu231*(-49);
assign relu2_weight43=bias2_relu20*(47)+bias2_relu21*(-18)+bias2_relu22*(30)+bias2_relu23*(-12)+bias2_relu24*(-13)+bias2_relu25*(-10)+bias2_relu26*(38)+bias2_relu27*(-11)+bias2_relu28*(-36)+bias2_relu29*(26)+bias2_relu210*(-17)+bias2_relu211*(27)+bias2_relu212*(38)+bias2_relu213*(32)+bias2_relu214*(-35)+bias2_relu215*(-28)+bias2_relu216*(-25)+bias2_relu217*(-20)+bias2_relu218*(-27)+bias2_relu219*(39)+bias2_relu220*(-47)+bias2_relu221*(-24)+bias2_relu222*(18)+bias2_relu223*(42)+bias2_relu224*(-3)+bias2_relu225*(-44)+bias2_relu226*(-11)+bias2_relu227*(24)+bias2_relu228*(-36)+bias2_relu229*(-55)+bias2_relu230*(-16)+bias2_relu231*(2);
assign relu2_weight44=bias2_relu20*(-53)+bias2_relu21*(-51)+bias2_relu22*(-72)+bias2_relu23*(-22)+bias2_relu24*(-6)+bias2_relu25*(17)+bias2_relu26*(-10)+bias2_relu27*(-39)+bias2_relu28*(-13)+bias2_relu29*(21)+bias2_relu210*(-32)+bias2_relu211*(26)+bias2_relu212*(-23)+bias2_relu213*(13)+bias2_relu214*(-79)+bias2_relu215*(43)+bias2_relu216*(51)+bias2_relu217*(53)+bias2_relu218*(47)+bias2_relu219*(-36)+bias2_relu220*(-3)+bias2_relu221*(-82)+bias2_relu222*(-22)+bias2_relu223*(23)+bias2_relu224*(0)+bias2_relu225*(24)+bias2_relu226*(-16)+bias2_relu227*(13)+bias2_relu228*(48)+bias2_relu229*(-13)+bias2_relu230*(-36)+bias2_relu231*(1);
assign relu2_weight45=bias2_relu20*(-32)+bias2_relu21*(32)+bias2_relu22*(25)+bias2_relu23*(-28)+bias2_relu24*(-17)+bias2_relu25*(31)+bias2_relu26*(17)+bias2_relu27*(-96)+bias2_relu28*(55)+bias2_relu29*(-65)+bias2_relu210*(-9)+bias2_relu211*(-17)+bias2_relu212*(0)+bias2_relu213*(5)+bias2_relu214*(2)+bias2_relu215*(-58)+bias2_relu216*(-71)+bias2_relu217*(-4)+bias2_relu218*(-15)+bias2_relu219*(33)+bias2_relu220*(-8)+bias2_relu221*(-11)+bias2_relu222*(41)+bias2_relu223*(-48)+bias2_relu224*(-6)+bias2_relu225*(-41)+bias2_relu226*(13)+bias2_relu227*(24)+bias2_relu228*(-20)+bias2_relu229*(51)+bias2_relu230*(18)+bias2_relu231*(24);
assign relu2_weight46=bias2_relu20*(24)+bias2_relu21*(19)+bias2_relu22*(-7)+bias2_relu23*(-16)+bias2_relu24*(30)+bias2_relu25*(-51)+bias2_relu26*(-42)+bias2_relu27*(-70)+bias2_relu28*(30)+bias2_relu29*(7)+bias2_relu210*(-27)+bias2_relu211*(-52)+bias2_relu212*(-77)+bias2_relu213*(36)+bias2_relu214*(-57)+bias2_relu215*(20)+bias2_relu216*(17)+bias2_relu217*(7)+bias2_relu218*(-14)+bias2_relu219*(25)+bias2_relu220*(-52)+bias2_relu221*(8)+bias2_relu222*(-49)+bias2_relu223*(12)+bias2_relu224*(-96)+bias2_relu225*(33)+bias2_relu226*(0)+bias2_relu227*(-81)+bias2_relu228*(37)+bias2_relu229*(45)+bias2_relu230*(44)+bias2_relu231*(-20);
assign relu2_weight47=bias2_relu20*(26)+bias2_relu21*(-12)+bias2_relu22*(-41)+bias2_relu23*(35)+bias2_relu24*(-42)+bias2_relu25*(6)+bias2_relu26*(-27)+bias2_relu27*(-24)+bias2_relu28*(1)+bias2_relu29*(7)+bias2_relu210*(19)+bias2_relu211*(64)+bias2_relu212*(-4)+bias2_relu213*(29)+bias2_relu214*(59)+bias2_relu215*(24)+bias2_relu216*(-3)+bias2_relu217*(-73)+bias2_relu218*(-9)+bias2_relu219*(-19)+bias2_relu220*(46)+bias2_relu221*(54)+bias2_relu222*(5)+bias2_relu223*(17)+bias2_relu224*(17)+bias2_relu225*(12)+bias2_relu226*(19)+bias2_relu227*(-43)+bias2_relu228*(-37)+bias2_relu229*(-15)+bias2_relu230*(-5)+bias2_relu231*(-41);
assign relu2_weight48=bias2_relu20*(-35)+bias2_relu21*(14)+bias2_relu22*(26)+bias2_relu23*(35)+bias2_relu24*(15)+bias2_relu25*(13)+bias2_relu26*(22)+bias2_relu27*(7)+bias2_relu28*(-13)+bias2_relu29*(37)+bias2_relu210*(1)+bias2_relu211*(-94)+bias2_relu212*(-15)+bias2_relu213*(9)+bias2_relu214*(7)+bias2_relu215*(-94)+bias2_relu216*(-87)+bias2_relu217*(37)+bias2_relu218*(-69)+bias2_relu219*(-46)+bias2_relu220*(-22)+bias2_relu221*(-49)+bias2_relu222*(-36)+bias2_relu223*(29)+bias2_relu224*(-21)+bias2_relu225*(2)+bias2_relu226*(-3)+bias2_relu227*(0)+bias2_relu228*(30)+bias2_relu229*(29)+bias2_relu230*(0)+bias2_relu231*(-27);
assign relu2_weight49=bias2_relu20*(4)+bias2_relu21*(-53)+bias2_relu22*(-7)+bias2_relu23*(22)+bias2_relu24*(-59)+bias2_relu25*(22)+bias2_relu26*(34)+bias2_relu27*(48)+bias2_relu28*(-45)+bias2_relu29*(-37)+bias2_relu210*(-122)+bias2_relu211*(-75)+bias2_relu212*(-30)+bias2_relu213*(-92)+bias2_relu214*(7)+bias2_relu215*(11)+bias2_relu216*(51)+bias2_relu217*(12)+bias2_relu218*(-1)+bias2_relu219*(-77)+bias2_relu220*(-3)+bias2_relu221*(-23)+bias2_relu222*(3)+bias2_relu223*(-12)+bias2_relu224*(31)+bias2_relu225*(-5)+bias2_relu226*(-17)+bias2_relu227*(17)+bias2_relu228*(2)+bias2_relu229*(-60)+bias2_relu230*(32)+bias2_relu231*(17);
wire [DATAWIDTH-1:0]   weight4_bias40;
wire [DATAWIDTH-1:0]   weight4_bias41;
wire [DATAWIDTH-1:0]   weight4_bias42;
wire [DATAWIDTH-1:0]   weight4_bias43;
wire [DATAWIDTH-1:0]   weight4_bias44;
wire [DATAWIDTH-1:0]   weight4_bias45;
wire [DATAWIDTH-1:0]   weight4_bias46;
wire [DATAWIDTH-1:0]   weight4_bias47;
wire [DATAWIDTH-1:0]   weight4_bias48;
wire [DATAWIDTH-1:0]   weight4_bias49;
assign weight4_bias40=relu2_weight40+(-11);
assign weight4_bias41=relu2_weight41+(9);
assign weight4_bias42=relu2_weight42+(-9);
assign weight4_bias43=relu2_weight43+(-7);
assign weight4_bias44=relu2_weight44+(29);
assign weight4_bias45=relu2_weight45+(32);
assign weight4_bias46=relu2_weight46+(-32);
assign weight4_bias47=relu2_weight47+(-15);
assign weight4_bias48=relu2_weight48+(-29);
assign weight4_bias49=relu2_weight49+(-2);
wire [4+DATAWIDTH-1:0] com_re01,com_re23,com_re45,com_re67,com_re89;
//check positive or negtive
assign com_re01=(result[0][DATAWIDTH-1]^result[1][DATAWIDTH-1]) ? 
                                                        ((result[0][DATAWIDTH-1]==1'b0)   ?   {4'd0,result[0]}:{4'd1,result[1]}):
                                                        ((result[0]>result[1]) ? {4'd0,result[0]}:{4'd1,result[1]});
assign com_re23=(result[2][DATAWIDTH-1]^result[3][DATAWIDTH-1]) ? 
                                                        ((result[2][DATAWIDTH-1]==1'b0)   ?   {4'd2,result[2]}:{4'd3,result[3]}):
                                                        ((result[2]>result[3]) ? {4'd2,result[2]}:{4'd3,result[3]});
assign com_re45=(result[4][DATAWIDTH-1]^result[5][DATAWIDTH-1]) ? 
                                                        ((result[4][DATAWIDTH-1]==1'b0)   ?   {4'd4,result[4]}:{4'd5,result[5]}):
                                                        ((result[4]>result[5]) ? {4'd4,result[4]}:{4'd5,result[5]});                                                        
assign com_re67=(result[6][DATAWIDTH-1]^result[7][DATAWIDTH-1]) ? 
                                                        ((result[6][DATAWIDTH-1]==1'b0)   ?   {4'd6,result[6]}:{4'd7,result[7]}):
                                                        ((result[6]>result[7]) ? {4'd6,result[6]}:{4'd7,result[7]});
assign com_re89=(result[8][DATAWIDTH-1]^result[9][DATAWIDTH-1]) ? 
                                                        ((result[8][DATAWIDTH-1]==1'b0)   ?   {4'd8,result[8]}:{4'd9,result[9]}):
                                                        ((result[8]>result[9]) ? {4'd8,result[8]}:{4'd9,result[9]});

wire [4+DATAWIDTH-1:0] com_re01_23,com_re45_67,com_re0123_4567,com_re01234567_89;
assign com_re01_23=(com_re01[DATAWIDTH-1]^com_re23[DATAWIDTH-1])   ?
                                                        ((com_re01[DATAWIDTH-1]==1'b0)  ?   com_re01:com_re23):
                                                        ((com_re01[DATAWIDTH-1:0]>com_re23[DATAWIDTH-1:0]) ?   com_re01:com_re23);
assign com_re45_67=(com_re45[DATAWIDTH-1]^com_re67[DATAWIDTH-1])   ?
                                                        ((com_re45[DATAWIDTH-1]==1'b0)  ?   com_re45:com_re67):
                                                        ((com_re45[DATAWIDTH-1:0]>com_re67[DATAWIDTH-1:0]) ?   com_re45:com_re67);
assign com_re0123_4567=(com_re01_23[DATAWIDTH-1]^com_re45_67[DATAWIDTH-1])   ?
                                                        ((com_re01_23[DATAWIDTH-1]==1'b0)  ?   com_re01_23:com_re45_67):
                                                        ((com_re01_23[DATAWIDTH-1:0]>com_re45_67[DATAWIDTH-1:0]) ?   com_re01_23:com_re45_67);
assign com_re01234567_89=(com_re0123_4567[DATAWIDTH-1]^com_re89[DATAWIDTH-1])   ?
                                                        ((com_re0123_4567[DATAWIDTH-1]==1'b0)  ?   com_re0123_4567:com_re89):
                                                        ((com_re0123_4567[DATAWIDTH-1:0]>com_re89[DATAWIDTH-1:0]) ?   com_re0123_4567:com_re89);


/////Eed Declatation////////
integer i;
always@(posedge clk or posedge rst)
   begin
       if(rst)
           begin
           for(i=0;i<784;i=i+1)
               begin
                   in_buf[i]<=0;
               end
           for(i=0;i<10;i=i+1)
               begin
                   result[i]<=0;
               end
               predict<=0;
           end
       else
       begin
           `include "in_buff.v"
            result[0]<=weight4_bias40;
            result[1]<=weight4_bias41;
            result[2]<=weight4_bias42;
            result[3]<=weight4_bias43;
            result[4]<=weight4_bias44;
            result[5]<=weight4_bias45;
            result[6]<=weight4_bias46;
            result[7]<=weight4_bias47;
            result[8]<=weight4_bias48;
            result[9]<=weight4_bias49;
           predict <=com_re01234567_89[4+DATAWIDTH-1:4+DATAWIDTH-1-3];       end
end


//wire declaration 

endmodule